magic
tech sky130A
timestamp 1731253424
<< metal1 >>
rect 11760 5125 11885 5130
rect 11760 5010 11765 5125
rect 11880 5010 11885 5125
rect 11760 5005 11885 5010
rect 11175 2715 11885 2840
rect 11175 510 11310 2715
rect 12655 2680 13090 2685
rect 12655 2565 12960 2680
rect 13085 2565 13090 2680
rect 12655 2560 13090 2565
rect 11760 1950 11885 1955
rect 11760 1835 11765 1950
rect 11880 1835 11885 1950
rect 11760 1830 11885 1835
rect 11175 380 15270 510
rect 15180 320 15270 380
rect 15180 270 15185 320
rect 15265 270 15270 320
rect 15180 265 15270 270
<< via1 >>
rect 11765 5010 11880 5125
rect 12960 2565 13085 2680
rect 11765 1835 11880 1950
rect 15185 270 15265 320
<< metal2 >>
rect 6762 19852 7454 19854
rect 6762 19823 7396 19852
rect 7449 19823 7454 19852
rect 6762 19822 7454 19823
rect 6762 18711 7740 18713
rect 6762 18682 7672 18711
rect 7725 18682 7740 18711
rect 6762 18681 7740 18682
rect 6762 17570 8006 17572
rect 6762 17541 7948 17570
rect 8001 17541 8006 17570
rect 6762 17540 8006 17541
rect 6762 16429 8282 16431
rect 6762 16400 8224 16429
rect 8277 16400 8282 16429
rect 6762 16399 8282 16400
rect 6762 15288 8558 15290
rect 6762 15259 8500 15288
rect 8553 15259 8558 15288
rect 6762 15258 8558 15259
rect 6762 14147 8834 14149
rect 6762 14118 8776 14147
rect 8829 14118 8834 14147
rect 6762 14117 8834 14118
rect 6762 13006 9110 13008
rect 6762 12977 9052 13006
rect 9105 12977 9110 13006
rect 6762 12976 9110 12977
rect 6762 11865 9386 11867
rect 6762 11836 9328 11865
rect 9381 11836 9386 11865
rect 6762 11835 9386 11836
rect 11635 5125 11885 5130
rect 11635 5010 11640 5125
rect 11755 5010 11765 5125
rect 11880 5010 11885 5125
rect 11635 5005 11885 5010
rect 12955 2680 13225 2685
rect 12955 2565 12960 2680
rect 13085 2565 13095 2680
rect 13220 2565 13225 2680
rect 12955 2560 13225 2565
rect 11635 1950 11885 1955
rect 11635 1835 11640 1950
rect 11755 1835 11765 1950
rect 11880 1835 11885 1950
rect 11635 1830 11885 1835
rect 15180 320 15270 325
rect 15180 270 15185 320
rect 15265 270 15270 320
rect 15180 245 15270 270
rect 15180 195 15185 245
rect 15265 195 15270 245
rect 15180 190 15270 195
<< via2 >>
rect 7396 19823 7449 19852
rect 7672 18682 7725 18711
rect 7948 17541 8001 17570
rect 8224 16400 8277 16429
rect 8500 15259 8553 15288
rect 8776 14118 8829 14147
rect 9052 12977 9105 13006
rect 9328 11836 9381 11865
rect 11640 5010 11755 5125
rect 13095 2565 13220 2680
rect 11640 1835 11755 1950
rect 15185 195 15265 245
<< metal3 >>
rect 7393 19858 7513 19861
rect 7393 19852 7477 19858
rect 7393 19823 7396 19852
rect 7449 19823 7477 19852
rect 7393 19818 7477 19823
rect 7510 19818 7513 19858
rect 7393 19816 7513 19818
rect 7669 18717 7789 18720
rect 7669 18711 7753 18717
rect 7669 18682 7672 18711
rect 7725 18682 7753 18711
rect 7669 18677 7753 18682
rect 7786 18677 7789 18717
rect 7669 18675 7789 18677
rect 7945 17576 8065 17579
rect 7945 17570 8029 17576
rect 7945 17541 7948 17570
rect 8001 17541 8029 17570
rect 7945 17536 8029 17541
rect 8062 17536 8065 17576
rect 7945 17534 8065 17536
rect 8221 16435 8341 16438
rect 8221 16429 8305 16435
rect 8221 16400 8224 16429
rect 8277 16400 8305 16429
rect 8221 16395 8305 16400
rect 8338 16395 8341 16435
rect 8221 16393 8341 16395
rect 8497 15294 8617 15297
rect 8497 15288 8581 15294
rect 8497 15259 8500 15288
rect 8553 15259 8581 15288
rect 8497 15254 8581 15259
rect 8614 15254 8617 15294
rect 8497 15252 8617 15254
rect 8773 14153 8893 14156
rect 8773 14147 8857 14153
rect 8773 14118 8776 14147
rect 8829 14118 8857 14147
rect 8773 14113 8857 14118
rect 8890 14113 8893 14153
rect 8773 14111 8893 14113
rect 9049 13012 9169 13015
rect 9049 13006 9133 13012
rect 9049 12977 9052 13006
rect 9105 12977 9133 13006
rect 9049 12972 9133 12977
rect 9166 12972 9169 13012
rect 9049 12970 9169 12972
rect 9325 11871 9445 11874
rect 9325 11865 9409 11871
rect 9325 11836 9328 11865
rect 9381 11836 9409 11865
rect 9325 11831 9409 11836
rect 9442 11831 9445 11871
rect 9325 11829 9445 11831
rect 100 5005 110 5130
rect 290 5125 11760 5130
rect 290 5010 11640 5125
rect 11755 5010 11760 5125
rect 290 5005 11760 5010
rect 13090 2680 13360 2685
rect 13090 2565 13095 2680
rect 13220 2565 13230 2680
rect 13355 2565 13360 2680
rect 13090 2560 13360 2565
rect 11510 1950 11760 1955
rect 11510 1835 11515 1950
rect 11630 1835 11640 1950
rect 11755 1835 11760 1950
rect 11510 1830 11760 1835
rect 15180 245 15270 250
rect 15180 195 15185 245
rect 15265 195 15270 245
rect 15180 170 15270 195
rect 15180 120 15185 170
rect 15265 120 15270 170
rect 15180 115 15270 120
<< via3 >>
rect 7477 19818 7510 19858
rect 7753 18677 7786 18717
rect 8029 17536 8062 17576
rect 8305 16395 8338 16435
rect 8581 15254 8614 15294
rect 8857 14113 8890 14153
rect 9133 12972 9166 13012
rect 9409 11831 9442 11871
rect 110 5005 290 5130
rect 13230 2565 13355 2680
rect 11515 1835 11630 1950
rect 15185 120 15265 170
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 100 5130 300 22076
rect 100 5005 110 5130
rect 290 5005 300 5130
rect 100 500 300 5005
rect 400 1955 600 22076
rect 7483 19861 7513 22576
rect 7474 19858 7513 19861
rect 7474 19818 7477 19858
rect 7510 19818 7513 19858
rect 7474 19816 7513 19818
rect 7759 18720 7789 22576
rect 7750 18717 7789 18720
rect 7750 18677 7753 18717
rect 7786 18677 7789 18717
rect 7750 18675 7789 18677
rect 8035 17579 8065 22576
rect 8026 17576 8065 17579
rect 8026 17536 8029 17576
rect 8062 17536 8065 17576
rect 8026 17534 8065 17536
rect 8311 16438 8341 22576
rect 8302 16435 8341 16438
rect 8302 16395 8305 16435
rect 8338 16395 8341 16435
rect 8302 16393 8341 16395
rect 8587 15297 8617 22576
rect 8578 15294 8617 15297
rect 8578 15254 8581 15294
rect 8614 15254 8617 15294
rect 8578 15252 8617 15254
rect 8863 14156 8893 22576
rect 8854 14153 8893 14156
rect 8854 14113 8857 14153
rect 8890 14113 8893 14153
rect 8854 14111 8893 14113
rect 9139 13015 9169 22576
rect 9130 13012 9169 13015
rect 9130 12972 9133 13012
rect 9166 12972 9169 13012
rect 9130 12970 9169 12972
rect 9415 11874 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22374 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 9406 11871 9445 11874
rect 9406 11831 9409 11871
rect 9442 11831 9445 11871
rect 9406 11829 9445 11831
rect 13225 2680 13360 2685
rect 13225 2565 13230 2680
rect 13355 2565 13360 2680
rect 400 1950 11635 1955
rect 400 1835 11515 1950
rect 11630 1835 11635 1950
rect 400 1830 11635 1835
rect 400 500 600 1830
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13225 0 13360 2565
rect 15180 170 15270 175
rect 15180 120 15185 170
rect 15265 120 15270 170
rect 15180 107 15270 120
rect 15178 0 15273 107
use input_stage  input_stage_0
timestamp 1731235174
transform 0 -1 9728 1 0 2180
box 46 160 1938 1275
use input_stage  input_stage_1
timestamp 1731235174
transform 0 -1 7787 1 0 2174
box 46 160 1938 1275
use inverter  inverter_0
timestamp 1728242959
transform 1 0 12080 0 1 1950
box -195 -120 615 3200
use tdc  tdc_0
timestamp 1730921041
transform 0 -1 6875 1 0 11141
box -6331 0 10295 3539
use variable_delay_dummy  variable_delay_dummy_0
timestamp 1731242716
transform 0 -1 8190 1 0 5543
box -3 0 3024 990
use variable_delay_short  variable_delay_short_0
timestamp 1731245751
transform 0 -1 12222 1 0 5729
box -3 0 8920 990
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 800 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
