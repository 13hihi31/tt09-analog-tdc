magic
tech sky130A
timestamp 1730652801
<< metal1 >>
rect 640 3323 1141 3371
rect 296 2785 352 2788
rect 296 2759 323 2785
rect 349 2759 352 2785
rect 296 2756 352 2759
rect 640 2628 1141 2676
<< via1 >>
rect 323 2759 349 2785
<< metal2 >>
rect 640 3277 1141 3309
rect 320 2785 352 2788
rect 320 2759 323 2785
rect 349 2759 352 2785
rect 320 2608 352 2759
rect 640 2692 1141 2724
rect 987 2608 1019 2692
rect 186 2576 352 2608
use delay_unit_2  delay_unit_2_0
timestamp 1730643297
transform 1 0 222 0 1 2699
box -222 -71 418 690
use saff_2  saff_2_0
timestamp 1730645859
transform 1 0 0 0 1 841
box 0 -841 1141 1767
<< end >>
