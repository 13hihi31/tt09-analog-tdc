magic
tech sky130A
magscale 1 2
timestamp 1731262231
<< metal1 >>
rect 9994 13290 10048 13300
rect 9990 13284 10052 13290
rect 9990 13214 9994 13284
rect 10048 13214 10052 13284
rect 9990 13208 10052 13214
rect 7804 10178 7858 10198
rect 15974 10196 16046 10202
rect 7800 10172 7862 10178
rect 7800 10102 7804 10172
rect 7858 10102 7862 10172
rect 7800 10096 7862 10102
rect 15148 10022 15516 10166
rect 15974 10134 15980 10196
rect 16042 10134 16046 10196
rect 15974 10128 16046 10134
rect 15148 8676 15292 10022
rect 15988 8572 16046 10128
rect 16342 8912 16408 10086
rect 16884 10038 17342 10182
rect 16342 8858 16348 8912
rect 16402 8858 16408 8912
rect 16342 8852 16408 8858
rect 17198 8676 17342 10038
rect 23646 9764 24088 9908
rect 24458 9894 24524 9900
rect 24458 9840 24464 9894
rect 24518 9840 24524 9894
rect 24458 9834 24524 9840
rect 23646 8678 23790 9764
rect 24480 8542 24524 9834
rect 25434 9816 25840 9960
rect 25696 8674 25840 9816
rect 16498 5570 16676 5576
rect 16498 5518 16502 5570
rect 16558 5518 16676 5570
rect 16498 5512 16676 5518
rect 16620 5292 16676 5512
rect 24378 5394 25174 5450
rect 25118 5262 25174 5394
rect 15814 4580 15916 4924
rect 15774 4562 16024 4580
rect 15774 4344 15790 4562
rect 16008 4344 16024 4562
rect 15774 4326 16024 4344
rect 16654 2472 16710 5108
rect 17240 3766 17342 4924
rect 24312 4580 24414 4896
rect 24272 4562 24522 4580
rect 24272 4344 24288 4562
rect 24506 4344 24522 4562
rect 24272 4326 24522 4344
rect 17152 3750 17402 3766
rect 17152 3528 17166 3750
rect 17386 3528 17402 3750
rect 17152 3516 17402 3528
rect 25152 2472 25208 5078
rect 25738 3766 25840 4932
rect 25648 3750 25898 3766
rect 25648 3528 25662 3750
rect 25882 3528 25898 3750
rect 25648 3516 25898 3528
rect 16654 2292 30540 2472
rect 30360 640 30540 2292
rect 30360 540 30370 640
rect 30530 540 30540 640
rect 30360 530 30540 540
<< via1 >>
rect 9994 13214 10048 13284
rect 7804 10102 7858 10172
rect 15980 10134 16042 10196
rect 16348 8858 16402 8912
rect 24464 9840 24518 9894
rect 16502 5518 16558 5570
rect 15790 4344 16008 4562
rect 24288 4344 24506 4562
rect 17166 3528 17386 3750
rect 25662 3528 25882 3750
rect 30370 540 30530 640
<< metal2 >>
rect 13524 39704 14908 39708
rect 13524 39646 14792 39704
rect 14898 39646 14908 39704
rect 13524 39644 14908 39646
rect 13524 37422 15480 37426
rect 13524 37364 15344 37422
rect 15450 37364 15480 37422
rect 13524 37362 15480 37364
rect 13524 35140 16012 35144
rect 13524 35082 15896 35140
rect 16002 35082 16012 35140
rect 13524 35080 16012 35082
rect 13524 32858 16564 32862
rect 13524 32800 16448 32858
rect 16554 32800 16564 32858
rect 13524 32798 16564 32800
rect 13524 30576 17116 30580
rect 13524 30518 17000 30576
rect 17106 30518 17116 30576
rect 13524 30516 17116 30518
rect 13524 28294 17668 28298
rect 13524 28236 17552 28294
rect 17658 28236 17668 28294
rect 13524 28234 17668 28236
rect 13524 26012 18220 26016
rect 13524 25954 18104 26012
rect 18210 25954 18220 26012
rect 13524 25952 18220 25954
rect 13524 23730 18772 23734
rect 13524 23672 18656 23730
rect 18762 23672 18772 23730
rect 13524 23670 18772 23672
rect 23298 21964 23702 21968
rect 23298 21906 23308 21964
rect 23414 21906 23702 21964
rect 23298 21904 23702 21906
rect 22746 18968 23702 18972
rect 22746 18910 22764 18968
rect 22870 18910 23702 18968
rect 22746 18908 23702 18910
rect 22354 16472 23704 16476
rect 22354 16414 22372 16472
rect 22478 16414 23704 16472
rect 22354 16412 23704 16414
rect 9990 13284 10052 13290
rect 9990 13214 9994 13284
rect 10048 13214 10052 13284
rect 7800 10172 7862 10178
rect 7800 10102 7804 10172
rect 7858 10102 7862 10172
rect 7800 8918 7862 10102
rect 9990 9277 10052 13214
rect 22154 13088 23692 13092
rect 22154 13030 22164 13088
rect 22270 13030 23692 13088
rect 22154 13028 23692 13030
rect 15964 10196 16046 10202
rect 15964 10134 15980 10196
rect 16042 10134 16046 10196
rect 15964 10102 16046 10134
rect 21992 10128 23690 10132
rect 21992 10070 22002 10128
rect 22108 10070 23690 10128
rect 21992 10068 23690 10070
rect 25129 9277 25195 9818
rect 9990 9211 25195 9277
rect 7800 8912 16408 8918
rect 7800 8858 16348 8912
rect 16402 8858 16408 8912
rect 7800 8852 16408 8858
rect 16586 8594 17594 8598
rect 16586 8536 17478 8594
rect 17584 8536 17594 8594
rect 16586 8534 17594 8536
rect 25084 8564 25948 8568
rect 25084 8506 25832 8564
rect 25938 8506 25948 8564
rect 25084 8504 25948 8506
rect 17084 8358 17874 8362
rect 17084 8300 17758 8358
rect 17864 8300 17874 8358
rect 17084 8298 17874 8300
rect 25582 8328 26500 8332
rect 25582 8270 26384 8328
rect 26490 8270 26500 8328
rect 25582 8268 26500 8270
rect 16586 7216 18152 7220
rect 16586 7158 18036 7216
rect 18142 7158 18152 7216
rect 16586 7156 18152 7158
rect 25084 7186 27052 7190
rect 25084 7128 26936 7186
rect 27042 7128 27052 7186
rect 25084 7126 27052 7128
rect 17084 6980 18496 6984
rect 17084 6922 18380 6980
rect 18486 6922 18496 6980
rect 17084 6920 18496 6922
rect 25582 6950 27604 6954
rect 25582 6892 27488 6950
rect 27594 6892 27604 6950
rect 25582 6890 27604 6892
rect 14760 5572 16562 5576
rect 14760 5514 14770 5572
rect 14876 5570 16562 5572
rect 14876 5518 16502 5570
rect 16558 5518 16562 5570
rect 14876 5514 16562 5518
rect 14760 5512 16562 5514
rect 15774 4562 16024 4580
rect 15774 4228 15790 4562
rect 16008 4228 16024 4562
rect 15774 4214 16024 4228
rect 24272 4562 24522 4580
rect 24272 4228 24288 4562
rect 24506 4228 24522 4562
rect 24272 4214 24522 4228
rect 17152 3750 17402 3766
rect 17152 3408 17166 3750
rect 17386 3408 17402 3750
rect 17152 3398 17402 3408
rect 25648 3750 25898 3766
rect 25648 3408 25662 3750
rect 25882 3408 25898 3750
rect 25648 3398 25898 3408
rect 30360 640 30540 650
rect 30360 540 30370 640
rect 30530 540 30540 640
rect 30360 490 30540 540
rect 30360 390 30370 490
rect 30530 390 30540 490
rect 30360 380 30540 390
<< via2 >>
rect 14792 39646 14898 39704
rect 15344 37364 15450 37422
rect 15896 35082 16002 35140
rect 16448 32800 16554 32858
rect 17000 30518 17106 30576
rect 17552 28236 17658 28294
rect 18104 25954 18210 26012
rect 18656 23672 18762 23730
rect 23308 21906 23414 21964
rect 22764 18910 22870 18968
rect 22372 16414 22478 16472
rect 22164 13030 22270 13088
rect 22002 10070 22108 10128
rect 17478 8536 17584 8594
rect 25832 8506 25938 8564
rect 17758 8300 17864 8358
rect 26384 8270 26490 8328
rect 18036 7158 18142 7216
rect 26936 7128 27042 7186
rect 18380 6922 18486 6980
rect 27488 6892 27594 6950
rect 14770 5514 14876 5572
rect 15790 4344 16008 4446
rect 15790 4228 16008 4344
rect 24288 4344 24506 4446
rect 24288 4228 24506 4344
rect 17166 3528 17386 3630
rect 17166 3408 17386 3528
rect 25662 3528 25882 3630
rect 25662 3408 25882 3528
rect 30370 390 30530 490
<< metal3 >>
rect 14786 39716 15026 39722
rect 14786 39704 14954 39716
rect 14786 39646 14792 39704
rect 14898 39646 14954 39704
rect 14786 39636 14954 39646
rect 15020 39636 15026 39716
rect 14786 39632 15026 39636
rect 15338 37434 15578 37440
rect 15338 37422 15506 37434
rect 15338 37364 15344 37422
rect 15450 37364 15506 37422
rect 15338 37354 15506 37364
rect 15572 37354 15578 37434
rect 15338 37350 15578 37354
rect 15890 35152 16130 35158
rect 15890 35140 16058 35152
rect 15890 35082 15896 35140
rect 16002 35082 16058 35140
rect 15890 35072 16058 35082
rect 16124 35072 16130 35152
rect 15890 35068 16130 35072
rect 16442 32870 16682 32876
rect 16442 32858 16610 32870
rect 16442 32800 16448 32858
rect 16554 32800 16610 32858
rect 16442 32790 16610 32800
rect 16676 32790 16682 32870
rect 16442 32786 16682 32790
rect 16994 30588 17234 30594
rect 16994 30576 17162 30588
rect 16994 30518 17000 30576
rect 17106 30518 17162 30576
rect 16994 30508 17162 30518
rect 17228 30508 17234 30588
rect 16994 30504 17234 30508
rect 17546 28306 17786 28312
rect 17546 28294 17714 28306
rect 17546 28236 17552 28294
rect 17658 28236 17714 28294
rect 17546 28226 17714 28236
rect 17780 28226 17786 28306
rect 17546 28222 17786 28226
rect 18098 26024 18338 26030
rect 18098 26012 18266 26024
rect 18098 25954 18104 26012
rect 18210 25954 18266 26012
rect 18098 25944 18266 25954
rect 18332 25944 18338 26024
rect 18098 25940 18338 25944
rect 18650 23742 18890 23748
rect 18650 23730 18818 23742
rect 18650 23672 18656 23730
rect 18762 23672 18818 23730
rect 18650 23662 18818 23672
rect 18884 23662 18890 23742
rect 18650 23658 18890 23662
rect 23180 21976 23420 21982
rect 23180 21896 23186 21976
rect 23252 21964 23420 21976
rect 23252 21906 23308 21964
rect 23414 21906 23420 21964
rect 23252 21896 23420 21906
rect 23180 21892 23420 21896
rect 22636 18980 22876 18986
rect 22636 18900 22642 18980
rect 22708 18968 22876 18980
rect 22708 18910 22764 18968
rect 22870 18910 22876 18968
rect 22708 18900 22876 18910
rect 22636 18896 22876 18900
rect 22244 16484 22484 16490
rect 22244 16404 22250 16484
rect 22316 16472 22484 16484
rect 22316 16414 22372 16472
rect 22478 16414 22484 16472
rect 22316 16404 22484 16414
rect 22244 16400 22484 16404
rect 22036 13100 22276 13106
rect 22036 13020 22042 13100
rect 22108 13088 22276 13100
rect 22108 13030 22164 13088
rect 22270 13030 22276 13088
rect 22108 13020 22276 13030
rect 22036 13016 22276 13020
rect 200 10010 220 10260
rect 580 10010 5808 10260
rect 21874 10140 22114 10146
rect 21874 10060 21880 10140
rect 21946 10128 22114 10140
rect 21946 10070 22002 10128
rect 22108 10070 22114 10128
rect 21946 10060 22114 10070
rect 21874 10056 22114 10060
rect 17472 8606 17712 8612
rect 17472 8594 17640 8606
rect 17472 8536 17478 8594
rect 17584 8536 17640 8594
rect 17472 8526 17640 8536
rect 17706 8526 17712 8606
rect 17472 8522 17712 8526
rect 25826 8576 26066 8582
rect 25826 8564 25994 8576
rect 25826 8506 25832 8564
rect 25938 8506 25994 8564
rect 25826 8496 25994 8506
rect 26060 8496 26066 8576
rect 25826 8492 26066 8496
rect 17752 8370 17992 8376
rect 17752 8358 17920 8370
rect 17752 8300 17758 8358
rect 17864 8300 17920 8358
rect 17752 8290 17920 8300
rect 17986 8290 17992 8370
rect 17752 8286 17992 8290
rect 26378 8340 26618 8346
rect 26378 8328 26546 8340
rect 26378 8270 26384 8328
rect 26490 8270 26546 8328
rect 26378 8260 26546 8270
rect 26612 8260 26618 8340
rect 26378 8256 26618 8260
rect 18030 7228 18270 7234
rect 18030 7216 18198 7228
rect 18030 7158 18036 7216
rect 18142 7158 18198 7216
rect 18030 7148 18198 7158
rect 18264 7148 18270 7228
rect 18030 7144 18270 7148
rect 26930 7198 27170 7204
rect 26930 7186 27098 7198
rect 26930 7128 26936 7186
rect 27042 7128 27098 7186
rect 26930 7118 27098 7128
rect 27164 7118 27170 7198
rect 26930 7114 27170 7118
rect 18374 6992 18614 6998
rect 18374 6980 18542 6992
rect 18374 6922 18380 6980
rect 18486 6922 18542 6980
rect 18374 6912 18542 6922
rect 18608 6912 18614 6992
rect 18374 6908 18614 6912
rect 27482 6962 27722 6968
rect 27482 6950 27650 6962
rect 27482 6892 27488 6950
rect 27594 6892 27650 6950
rect 27482 6882 27650 6892
rect 27716 6882 27722 6962
rect 27482 6878 27722 6882
rect 14642 5584 14882 5590
rect 14642 5504 14648 5584
rect 14714 5572 14882 5584
rect 14714 5514 14770 5572
rect 14876 5514 14882 5572
rect 14714 5504 14882 5514
rect 14642 5500 14882 5504
rect 198 4214 220 4464
rect 580 4446 24522 4464
rect 580 4228 15790 4446
rect 16008 4228 24288 4446
rect 24506 4228 24522 4446
rect 580 4214 24522 4228
rect 17152 3636 17402 3648
rect 25648 3636 25898 3648
rect 17151 3630 17402 3636
rect 17151 3300 17166 3630
rect 17386 3300 17402 3630
rect 17151 3290 17402 3300
rect 25647 3630 25898 3636
rect 25647 3300 25662 3630
rect 25882 3300 25898 3630
rect 25647 3290 25898 3300
rect 30360 490 30540 500
rect 30360 390 30370 490
rect 30530 390 30540 490
rect 30360 340 30540 390
rect 30360 240 30370 340
rect 30530 240 30540 340
rect 30360 230 30540 240
<< via3 >>
rect 14954 39636 15020 39716
rect 15506 37354 15572 37434
rect 16058 35072 16124 35152
rect 16610 32790 16676 32870
rect 17162 30508 17228 30588
rect 17714 28226 17780 28306
rect 18266 25944 18332 26024
rect 18818 23662 18884 23742
rect 23186 21896 23252 21976
rect 22642 18900 22708 18980
rect 22250 16404 22316 16484
rect 22042 13020 22108 13100
rect 220 10010 580 10260
rect 21880 10060 21946 10140
rect 17640 8526 17706 8606
rect 25994 8496 26060 8576
rect 17920 8290 17986 8370
rect 26546 8260 26612 8340
rect 18198 7148 18264 7228
rect 27098 7118 27164 7198
rect 18542 6912 18608 6992
rect 27650 6882 27716 6962
rect 14648 5504 14714 5584
rect 220 4214 580 4464
rect 17166 3408 17386 3526
rect 17166 3300 17386 3408
rect 25662 3408 25882 3526
rect 25662 3300 25882 3408
rect 30370 240 30530 340
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 200 10260 600 44152
rect 200 10010 220 10260
rect 580 10010 600 10260
rect 200 4464 600 10010
rect 200 4214 220 4464
rect 580 4214 600 4464
rect 200 1000 600 4214
rect 800 3540 1200 44152
rect 14966 39722 15026 45152
rect 14948 39716 15026 39722
rect 14948 39636 14954 39716
rect 15020 39636 15026 39716
rect 14948 39632 15026 39636
rect 15518 37440 15578 45152
rect 15500 37434 15578 37440
rect 15500 37354 15506 37434
rect 15572 37354 15578 37434
rect 15500 37350 15578 37354
rect 16070 35158 16130 45152
rect 16052 35152 16130 35158
rect 16052 35072 16058 35152
rect 16124 35072 16130 35152
rect 16052 35068 16130 35072
rect 16622 32876 16682 45152
rect 16604 32870 16682 32876
rect 16604 32790 16610 32870
rect 16676 32790 16682 32870
rect 16604 32786 16682 32790
rect 17174 30594 17234 45152
rect 17156 30588 17234 30594
rect 17156 30508 17162 30588
rect 17228 30508 17234 30588
rect 17156 30504 17234 30508
rect 17726 28312 17786 45152
rect 17708 28306 17786 28312
rect 17708 28226 17714 28306
rect 17780 28226 17786 28306
rect 17708 28222 17786 28226
rect 18278 26030 18338 45152
rect 18260 26024 18338 26030
rect 18260 25944 18266 26024
rect 18332 25944 18338 26024
rect 18260 25940 18338 25944
rect 18830 23748 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 32176 20546 45152
rect 18812 23742 18890 23748
rect 18812 23662 18818 23742
rect 18884 23662 18890 23742
rect 18812 23658 18890 23662
rect 20122 32116 20546 32176
rect 20122 13260 20182 32116
rect 21038 31746 21098 45152
rect 17356 13200 20182 13260
rect 20490 31686 21098 31746
rect 17356 9688 17416 13200
rect 20490 12952 20550 31686
rect 21590 31308 21650 45152
rect 14642 9628 17416 9688
rect 17652 12892 20550 12952
rect 20798 31248 21650 31308
rect 14642 5590 14702 9628
rect 17652 8612 17712 12892
rect 20798 12686 20858 31248
rect 22142 30932 22202 45152
rect 17634 8606 17712 8612
rect 17634 8526 17640 8606
rect 17706 8526 17712 8606
rect 17634 8522 17712 8526
rect 17932 12626 20858 12686
rect 21188 30872 22202 30932
rect 17932 8376 17992 12626
rect 21188 12394 21248 30872
rect 22694 30470 22754 45152
rect 17914 8370 17992 8376
rect 17914 8290 17920 8370
rect 17986 8290 17992 8370
rect 17914 8286 17992 8290
rect 18210 12334 21248 12394
rect 21479 30410 22754 30470
rect 18210 7234 18270 12334
rect 21479 12041 21540 30410
rect 23246 29882 23306 45152
rect 18192 7228 18270 7234
rect 18192 7148 18198 7228
rect 18264 7148 18270 7228
rect 18192 7144 18270 7148
rect 18554 11980 21540 12041
rect 21874 29822 23306 29882
rect 18554 7018 18615 11980
rect 21874 10146 21934 29822
rect 23798 29616 23858 45152
rect 22036 29556 23858 29616
rect 22036 13106 22096 29556
rect 24350 29386 24410 45152
rect 22244 29326 24410 29386
rect 22244 16490 22304 29326
rect 24902 29066 24962 45152
rect 22636 29006 24962 29066
rect 22636 18986 22696 29006
rect 25454 28658 25514 45152
rect 23180 28598 25514 28658
rect 23180 21982 23240 28598
rect 23180 21976 23258 21982
rect 23180 21896 23186 21976
rect 23252 21896 23258 21976
rect 23180 21892 23258 21896
rect 22636 18980 22714 18986
rect 22636 18900 22642 18980
rect 22708 18900 22714 18980
rect 22636 18896 22714 18900
rect 22244 16484 22322 16490
rect 22244 16404 22250 16484
rect 22316 16404 22322 16484
rect 22244 16400 22322 16404
rect 22036 13100 22114 13106
rect 22036 13020 22042 13100
rect 22108 13020 22114 13100
rect 22036 13016 22114 13020
rect 21874 10140 21952 10146
rect 21874 10060 21880 10140
rect 21946 10060 21952 10140
rect 21874 10056 21952 10060
rect 26006 8582 26066 45152
rect 25988 8576 26066 8582
rect 25988 8496 25994 8576
rect 26060 8496 26066 8576
rect 25988 8492 26066 8496
rect 26558 8346 26618 45152
rect 26540 8340 26618 8346
rect 26540 8260 26546 8340
rect 26612 8260 26618 8340
rect 26540 8256 26618 8260
rect 27110 7204 27170 45152
rect 27092 7198 27170 7204
rect 27092 7118 27098 7198
rect 27164 7118 27170 7198
rect 27092 7114 27170 7118
rect 18554 6998 18614 7018
rect 18536 6992 18614 6998
rect 18536 6912 18542 6992
rect 18608 6912 18614 6992
rect 27662 6968 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 18536 6908 18614 6912
rect 27644 6962 27722 6968
rect 27644 6882 27650 6962
rect 27716 6882 27722 6962
rect 27644 6878 27722 6882
rect 14642 5584 14720 5590
rect 14642 5504 14648 5584
rect 14714 5504 14720 5584
rect 14642 5500 14720 5504
rect 800 3526 25898 3540
rect 800 3300 17166 3526
rect 17386 3300 25662 3526
rect 25882 3300 25898 3526
rect 800 3290 25898 3300
rect 800 1000 1200 3290
rect 30360 340 30540 350
rect 30360 240 30370 340
rect 30530 240 30540 340
rect 30360 214 30540 240
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30356 0 30546 214
use input_stage  input_stage_0
timestamp 1731235174
transform 0 -1 17662 1 0 4832
box 92 320 3876 2550
use input_stage  input_stage_1
timestamp 1731235174
transform 0 -1 26160 1 0 4802
box 92 320 3876 2550
use tdc  tdc_0
timestamp 1730921041
transform 0 -1 13750 1 0 22282
box -12662 0 20590 7078
use variable_delay_dummy  variable_delay_dummy_0
timestamp 1731242716
transform 0 -1 17052 1 0 10020
box -6 0 6048 1980
use variable_delay_short  variable_delay_short_0
timestamp 1731245751
transform 0 -1 25612 1 0 9752
box -6 0 17840 1980
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
