magic
tech sky130A
magscale 1 2
timestamp 1730537487
<< nwell >>
rect 5844 -388 7140 -152
rect 5844 -1112 5990 -388
rect 6442 -1112 6660 -388
rect 6996 -1112 7140 -388
<< pwell >>
rect 5844 -1780 7140 -1112
<< psubdiff >>
rect 5918 -1254 5954 -1230
rect 6472 -1162 6508 -1138
rect 7032 -1254 7068 -1230
rect 5886 -1780 5910 -1678
rect 7076 -1780 7100 -1678
<< nsubdiff >>
rect 5880 -304 5904 -202
rect 7080 -304 7104 -202
rect 5918 -448 5954 -304
rect 5918 -1076 5954 -1052
rect 6472 -448 6508 -304
rect 6472 -1076 6508 -1052
rect 7032 -448 7068 -304
rect 7032 -1076 7068 -1052
<< psubdiffcont >>
rect 5918 -1678 5954 -1254
rect 6472 -1678 6508 -1162
rect 7032 -1678 7068 -1254
rect 5910 -1780 7076 -1678
<< nsubdiffcont >>
rect 5904 -304 7080 -202
rect 5918 -1052 5954 -448
rect 6472 -1052 6508 -448
rect 7032 -1052 7068 -448
<< poly >>
rect 6226 -356 6292 -340
rect 6226 -390 6242 -356
rect 6276 -390 6292 -356
rect 6226 -406 6292 -390
rect 6242 -426 6272 -406
rect 6688 -354 6754 -338
rect 6688 -388 6704 -354
rect 6738 -388 6754 -354
rect 6688 -404 6754 -388
rect 6708 -424 6738 -404
rect 5966 -1096 6096 -1066
rect 5966 -1132 5996 -1096
rect 5900 -1148 5996 -1132
rect 6154 -1138 6184 -1076
rect 5900 -1182 5916 -1148
rect 5950 -1182 5996 -1148
rect 5900 -1198 5996 -1182
rect 6088 -1150 6184 -1138
rect 6088 -1184 6104 -1150
rect 6138 -1166 6184 -1150
rect 6330 -1090 6360 -1076
rect 6330 -1102 6396 -1090
rect 6330 -1136 6346 -1102
rect 6380 -1136 6396 -1102
rect 6330 -1148 6396 -1136
rect 6138 -1184 6272 -1166
rect 6088 -1196 6272 -1184
rect 5966 -1238 5996 -1198
rect 5966 -1268 6096 -1238
rect 6242 -1258 6272 -1196
rect 6330 -1258 6360 -1148
rect 6154 -1554 6184 -1508
rect 6004 -1570 6184 -1554
rect 6004 -1604 6020 -1570
rect 6054 -1584 6184 -1570
rect 6054 -1604 6070 -1584
rect 6004 -1620 6070 -1604
rect 6620 -1194 6650 -1076
rect 6796 -1138 6826 -1076
rect 6884 -1096 7014 -1066
rect 6984 -1132 7014 -1096
rect 6796 -1150 6892 -1138
rect 6796 -1166 6842 -1150
rect 6584 -1206 6650 -1194
rect 6584 -1240 6600 -1206
rect 6634 -1240 6650 -1206
rect 6584 -1252 6650 -1240
rect 6620 -1260 6650 -1252
rect 6708 -1184 6842 -1166
rect 6876 -1184 6892 -1150
rect 6708 -1196 6892 -1184
rect 6984 -1148 7080 -1132
rect 6984 -1182 7030 -1148
rect 7064 -1182 7080 -1148
rect 6708 -1258 6738 -1196
rect 6984 -1198 7080 -1182
rect 6984 -1238 7014 -1198
rect 6884 -1268 7014 -1238
rect 6796 -1556 6826 -1510
rect 6796 -1572 6976 -1556
rect 6796 -1586 6926 -1572
rect 6910 -1606 6926 -1586
rect 6960 -1606 6976 -1572
rect 6910 -1622 6976 -1606
<< polycont >>
rect 6242 -390 6276 -356
rect 6704 -388 6738 -354
rect 5916 -1182 5950 -1148
rect 6104 -1184 6138 -1150
rect 6346 -1136 6380 -1102
rect 6020 -1604 6054 -1570
rect 6600 -1240 6634 -1206
rect 6842 -1184 6876 -1150
rect 7030 -1182 7064 -1148
rect 6926 -1606 6960 -1572
<< locali >>
rect 5880 -304 5904 -202
rect 7080 -304 7104 -202
rect 5918 -448 5954 -304
rect 6226 -356 6292 -350
rect 6226 -390 6242 -356
rect 6276 -390 6292 -356
rect 6226 -396 6292 -390
rect 5918 -1076 5954 -1052
rect 6472 -448 6508 -304
rect 6688 -354 6754 -348
rect 6688 -388 6704 -354
rect 6738 -388 6754 -354
rect 6688 -394 6754 -388
rect 6472 -1076 6508 -1052
rect 7032 -448 7068 -304
rect 7032 -1076 7068 -1052
rect 6330 -1102 6396 -1096
rect 6330 -1136 6346 -1102
rect 6380 -1136 6396 -1102
rect 6330 -1142 6396 -1136
rect 5900 -1148 5966 -1142
rect 5900 -1182 5916 -1148
rect 5950 -1182 5966 -1148
rect 5900 -1188 5966 -1182
rect 6088 -1150 6154 -1146
rect 6088 -1184 6104 -1150
rect 6138 -1184 6154 -1150
rect 6088 -1188 6154 -1184
rect 6472 -1162 6508 -1138
rect 5918 -1254 5954 -1230
rect 6826 -1150 6892 -1144
rect 6826 -1184 6842 -1150
rect 6876 -1184 6892 -1150
rect 6826 -1190 6892 -1184
rect 7014 -1148 7080 -1142
rect 7014 -1182 7030 -1148
rect 7064 -1182 7080 -1148
rect 7014 -1188 7080 -1182
rect 6584 -1206 6650 -1200
rect 6584 -1240 6600 -1206
rect 6634 -1240 6650 -1206
rect 6584 -1246 6650 -1240
rect 6004 -1570 6070 -1564
rect 6004 -1604 6020 -1570
rect 6054 -1604 6070 -1570
rect 6004 -1610 6070 -1604
rect 7032 -1254 7068 -1230
rect 6910 -1572 6976 -1566
rect 6910 -1606 6926 -1572
rect 6960 -1606 6976 -1572
rect 6910 -1612 6976 -1606
rect 5886 -1780 5910 -1678
rect 7076 -1780 7100 -1678
<< viali >>
rect 5904 -298 7080 -208
rect 6242 -390 6276 -356
rect 5918 -1052 5954 -448
rect 6704 -388 6738 -354
rect 6472 -1052 6508 -448
rect 7032 -1052 7068 -448
rect 6346 -1136 6380 -1102
rect 5916 -1182 5950 -1148
rect 6104 -1184 6138 -1150
rect 5918 -1648 5954 -1322
rect 6842 -1184 6876 -1150
rect 7030 -1182 7064 -1148
rect 6600 -1240 6634 -1206
rect 6020 -1604 6054 -1570
rect 6472 -1648 6508 -1300
rect 6926 -1606 6960 -1572
rect 7032 -1648 7068 -1322
rect 5910 -1772 7076 -1686
<< metal1 >>
rect 5844 -208 7140 -202
rect 5844 -298 5904 -208
rect 7080 -298 7140 -208
rect 5844 -304 7140 -298
rect 5912 -448 5960 -304
rect 5994 -346 6060 -340
rect 5994 -400 6000 -346
rect 6054 -400 6060 -346
rect 5994 -406 6060 -400
rect 5912 -1052 5918 -448
rect 5954 -1052 5960 -448
rect 6014 -450 6060 -406
rect 6102 -450 6148 -304
rect 6226 -346 6292 -340
rect 6226 -400 6232 -346
rect 6286 -400 6292 -346
rect 6226 -406 6292 -400
rect 6366 -450 6412 -304
rect 6466 -448 6514 -304
rect 5912 -1064 5960 -1052
rect 5900 -1138 5966 -1132
rect 5900 -1192 5906 -1138
rect 5960 -1192 5966 -1138
rect 5900 -1198 5966 -1192
rect 6014 -1284 6060 -1050
rect 6088 -1140 6154 -1134
rect 6088 -1194 6094 -1140
rect 6148 -1194 6154 -1140
rect 6088 -1200 6154 -1194
rect 6190 -1200 6236 -1050
rect 6466 -1052 6472 -448
rect 6508 -1052 6514 -448
rect 6568 -450 6614 -304
rect 6688 -344 6754 -338
rect 6688 -398 6694 -344
rect 6748 -398 6754 -344
rect 6688 -404 6754 -398
rect 6832 -450 6878 -304
rect 6920 -344 6986 -338
rect 6920 -398 6926 -344
rect 6980 -398 6986 -344
rect 6920 -404 6986 -398
rect 6920 -450 6966 -404
rect 7026 -448 7074 -304
rect 6466 -1064 6514 -1052
rect 6744 -1096 6790 -1050
rect 6330 -1102 6790 -1096
rect 6330 -1136 6346 -1102
rect 6380 -1136 6790 -1102
rect 6330 -1142 6790 -1136
rect 6190 -1206 6650 -1200
rect 6190 -1240 6600 -1206
rect 6634 -1240 6650 -1206
rect 6190 -1246 6650 -1240
rect 6190 -1284 6236 -1246
rect 6744 -1284 6790 -1142
rect 6826 -1140 6892 -1134
rect 6826 -1194 6832 -1140
rect 6886 -1194 6892 -1140
rect 6826 -1200 6892 -1194
rect 6920 -1284 6966 -1050
rect 7026 -1052 7032 -448
rect 7068 -1052 7074 -448
rect 7026 -1064 7074 -1052
rect 7014 -1138 7080 -1132
rect 7014 -1192 7020 -1138
rect 7074 -1192 7080 -1138
rect 7014 -1198 7080 -1192
rect 6466 -1300 6514 -1284
rect 5912 -1322 5960 -1310
rect 5912 -1648 5918 -1322
rect 5954 -1648 5960 -1322
rect 6014 -1570 6060 -1484
rect 6014 -1604 6020 -1570
rect 6054 -1604 6060 -1570
rect 6014 -1620 6060 -1604
rect 5912 -1678 5960 -1648
rect 6102 -1678 6148 -1484
rect 6190 -1554 6236 -1484
rect 6190 -1560 6254 -1554
rect 6190 -1612 6196 -1560
rect 6248 -1612 6254 -1560
rect 6190 -1618 6254 -1612
rect 6366 -1678 6412 -1484
rect 6466 -1648 6472 -1300
rect 6508 -1648 6514 -1300
rect 7026 -1322 7074 -1310
rect 6466 -1678 6514 -1648
rect 6568 -1678 6614 -1484
rect 6744 -1556 6790 -1484
rect 6726 -1562 6790 -1556
rect 6726 -1614 6732 -1562
rect 6784 -1614 6790 -1562
rect 6726 -1620 6790 -1614
rect 6832 -1678 6878 -1484
rect 6920 -1572 6966 -1484
rect 6920 -1606 6926 -1572
rect 6960 -1606 6966 -1572
rect 6920 -1622 6966 -1606
rect 7026 -1648 7032 -1322
rect 7068 -1648 7074 -1322
rect 7026 -1678 7074 -1648
rect 5844 -1686 7140 -1678
rect 5844 -1772 5910 -1686
rect 7076 -1772 7140 -1686
rect 5844 -1780 7140 -1772
<< via1 >>
rect 6000 -400 6054 -346
rect 6232 -356 6286 -346
rect 6232 -390 6242 -356
rect 6242 -390 6276 -356
rect 6276 -390 6286 -356
rect 6232 -400 6286 -390
rect 5906 -1148 5960 -1138
rect 5906 -1182 5916 -1148
rect 5916 -1182 5950 -1148
rect 5950 -1182 5960 -1148
rect 5906 -1192 5960 -1182
rect 6094 -1150 6148 -1140
rect 6094 -1184 6104 -1150
rect 6104 -1184 6138 -1150
rect 6138 -1184 6148 -1150
rect 6094 -1194 6148 -1184
rect 6694 -354 6748 -344
rect 6694 -388 6704 -354
rect 6704 -388 6738 -354
rect 6738 -388 6748 -354
rect 6694 -398 6748 -388
rect 6926 -398 6980 -344
rect 6832 -1150 6886 -1140
rect 6832 -1184 6842 -1150
rect 6842 -1184 6876 -1150
rect 6876 -1184 6886 -1150
rect 6832 -1194 6886 -1184
rect 7020 -1148 7074 -1138
rect 7020 -1182 7030 -1148
rect 7030 -1182 7064 -1148
rect 7064 -1182 7074 -1148
rect 7020 -1192 7074 -1182
rect 6196 -1612 6248 -1560
rect 6732 -1614 6784 -1562
<< metal2 >>
rect 5844 -1132 5890 -324
rect 5994 -346 6292 -340
rect 5994 -400 6000 -346
rect 6054 -400 6232 -346
rect 6286 -400 6292 -346
rect 6688 -344 6986 -338
rect 5994 -406 6292 -400
rect 5844 -1138 5966 -1132
rect 5844 -1178 5906 -1138
rect 5900 -1192 5906 -1178
rect 5960 -1192 5966 -1138
rect 5900 -1198 5966 -1192
rect 6088 -1140 6154 -1134
rect 6088 -1194 6094 -1140
rect 6148 -1146 6154 -1140
rect 6416 -1146 6462 -360
rect 6148 -1194 6462 -1146
rect 6518 -1148 6564 -360
rect 6688 -398 6694 -344
rect 6748 -398 6926 -344
rect 6980 -398 6986 -344
rect 6688 -404 6986 -398
rect 7094 -1132 7140 -332
rect 6826 -1140 6892 -1134
rect 6826 -1148 6832 -1140
rect 6518 -1194 6832 -1148
rect 6886 -1194 6892 -1140
rect 6088 -1200 6154 -1194
rect 6826 -1200 6892 -1194
rect 7014 -1138 7140 -1132
rect 7014 -1192 7020 -1138
rect 7074 -1178 7140 -1138
rect 7074 -1192 7080 -1178
rect 7014 -1198 7080 -1192
rect 6190 -1560 6254 -1554
rect 6190 -1612 6196 -1560
rect 6248 -1612 6254 -1560
rect 6190 -1618 6254 -1612
rect 6726 -1562 6790 -1556
rect 6726 -1614 6732 -1562
rect 6784 -1614 6790 -1562
rect 6726 -1620 6790 -1614
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1730191042
transform 1 0 6081 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1730191042
transform 1 0 6169 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1730191042
transform 1 0 6257 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1730191042
transform 1 0 6345 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1730191042
transform 1 0 6635 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1730191042
transform 1 0 6723 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_6
timestamp 1730191042
transform 1 0 6811 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_7
timestamp 1730191042
transform 1 0 6899 0 1 -1384
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_0
timestamp 1730191042
transform 1 0 6081 0 1 -750
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_1
timestamp 1730191042
transform 1 0 6169 0 1 -750
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_2
timestamp 1730191042
transform 1 0 6257 0 1 -750
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_3
timestamp 1730191042
transform 1 0 6345 0 1 -750
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_4
timestamp 1730191042
transform 1 0 6635 0 1 -750
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_5
timestamp 1730191042
transform 1 0 6723 0 1 -750
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_6
timestamp 1730191042
transform 1 0 6811 0 1 -750
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_7
timestamp 1730191042
transform 1 0 6899 0 1 -750
box -109 -362 109 362
<< labels >>
rlabel metal2 6416 -408 6462 -360 0 a1
port 1 nsew
rlabel metal2 6518 -408 6564 -360 0 b1
port 3 nsew
rlabel metal2 6190 -1618 6254 -1554 0 c
port 5 nsew
rlabel metal2 6726 -1620 6790 -1556 0 nc
port 6 nsew
rlabel metal1 5844 -238 5880 -202 0 VDD
port 7 nsew
rlabel metal1 5844 -1720 5886 -1678 0 VSS
port 8 nsew
rlabel metal2 7094 -380 7140 -332 0 a2
port 2 nsew
rlabel metal2 5844 -372 5890 -324 0 b2
port 4 nsew
<< end >>
