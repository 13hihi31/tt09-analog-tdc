magic
tech sky130A
timestamp 1730838452
<< metal1 >>
rect -4829 3323 -4688 3371
rect -208 3323 -45 3371
rect -5353 3289 -5318 3292
rect -5353 3260 -5350 3289
rect -5321 3260 -5318 3289
rect -5353 3257 -5318 3260
rect -4874 2676 -4829 2748
rect -4874 2628 -4688 2676
rect -4874 1701 -4829 2628
rect -382 2228 -29 2276
rect -4874 1653 -4496 1701
rect -427 51 -382 1653
rect -427 0 150 51
<< via1 >>
rect -5350 3260 -5321 3289
rect 75 2512 117 2555
<< metal2 >>
rect -5353 3428 -4726 3464
rect -5353 3289 -5318 3428
rect -5353 3260 -5350 3289
rect -5321 3260 -5318 3289
rect -4762 3309 -4726 3428
rect -4762 3277 -4688 3309
rect -208 3277 256 3309
rect -5353 3257 -5318 3260
rect -4883 2827 -4688 2862
rect -140 2772 256 2804
rect -140 2724 -108 2772
rect -208 2692 -108 2724
rect -233 2555 121 2558
rect -233 2512 75 2555
rect 117 2512 121 2555
rect -233 2508 121 2512
rect -233 1785 -183 2508
rect -471 1732 -183 1785
use diff_gen  diff_gen_0
timestamp 1730821783
transform 1 0 -4688 0 1 2628
box 0 0 4480 761
use start_buffer  start_buffer_0
timestamp 1730835638
transform 1 0 -6043 0 1 2748
box 0 0 1214 641
use stop_buffer  stop_buffer_0
timestamp 1730753331
transform 1 0 -4496 0 1 1653
box 0 0 4114 641
use vernier_delay_line  vernier_delay_line_0
timestamp 1730836525
transform 1 0 256 0 1 0
box -301 0 9768 3389
<< end >>
