* NGSPICE file created from tt_um_13hihi31_tdc_parax.ext - technology: sky130A

.subckt tt_um_13hihi31_tdc_parax clk ena rst_n ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[1]
+ ui_in[5] uo_out[7] ui_in[7] uio_in[0] uo_out[6] ui_in[4] uo_out[5] ui_in[0] uo_out[4]
+ uo_out[0] ui_in[3] uo_out[3] ui_in[6] ui_in[2] VGND VDPWR ui_in[1] uo_out[2] ua[0]
X0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 VDPWR.t460 VDPWR.t459 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1 tdc_0.start_buffer_0.start_delay.t6 tdc_0.start_buffer_0.start_buff.t10 VDPWR.t89 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X2 a_24240_14314# variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t2 VDPWR.t503 VDPWR.t502 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X3 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 VGND.t24 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X4 tdc_0.vernier_delay_line_0.stop_strong.t15 a_9330_16954.t8 VGND.t250 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5 a_10958_39338.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 a_10108_39954.t4 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X6 a_10108_28544.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X7 VDPWR.t241 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12420_30598# VDPWR.t240 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X8 VGND.t416 input_stage_1.fine_delay_unit_0.in a_24790_6936# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X9 a_10958_23364.t6 tdc_0.vernier_delay_line_0.stop_strong.t32 VGND.t301 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X10 a_24240_11366# variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t2 VDPWR.t340 VDPWR.t339 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 a_13254_26412# VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X12 tdc_0.vernier_delay_line_0.stop_strong.t31 a_9330_16954.t9 VDPWR.t107 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X13 a_10108_35390.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 a_13254_35540# VGND.t306 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X15 VDPWR.t199 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 VDPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X16 VGND.t86 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t2 a_25060_21092# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X17 a_10108_39426# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 a_10958_39338.t12 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X18 VDPWR.t352 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t2 a_24240_26106# VDPWR.t351 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X19 a_10958_37056.t10 tdc_0.vernier_delay_line_0.stop_strong.t33 VGND.t155 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X20 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 a_10108_26262.t5 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X21 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t1 VDPWR.t451 VDPWR.t452 VDPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X22 VGND.t156 tdc_0.vernier_delay_line_0.stop_strong.t34 a_10958_23364.t5 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X23 a_9330_14344# a_9330_14054# VGND.t187 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X24 uo_out[6].t3 a_12310_37398# VGND.t186 VGND.t185 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X25 VGND.t230 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VGND.t229 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X26 a_25060_24040# variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t2 VGND.t358 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X27 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 a_10108_35390.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X28 a_9330_16954.t3 a_9330_15794# VGND.t540 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X29 VDPWR.t413 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t3 a_24240_23158# VDPWR.t412 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X30 a_7140_10670# variable_delay_dummy_0.out VDPWR.t568 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X31 variable_delay_short_0.in a_23820_8460# VGND.t81 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X32 a_25060_21092# variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t3 VGND.t87 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X33 VGND.t490 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X34 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t7 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t8 VDPWR.t179 VDPWR.t178 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X35 VDPWR.t312 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t8 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t1 VDPWR.t311 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X36 a_10108_39426# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 a_10958_39338.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X37 a_10958_37056.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 a_10108_37144# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X38 VGND.t168 tdc_0.vernier_delay_line_0.stop_strong.t35 a_10958_34774.t9 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X39 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t7 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t8 VDPWR.t545 VDPWR.t544 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X40 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12308_33296# a_12420_33258# VDPWR.t476 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X41 VGND.t415 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 VGND.t414 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X42 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 VGND.t51 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X43 a_13254_35162# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 uo_out[5].t1 VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X44 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 VDPWR.t378 VDPWR.t377 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X45 a_25060_18144# variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t2 VGND.t541 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X46 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t0 ui_in[5].t0 VDPWR.t184 VDPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X47 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t5 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t8 VDPWR.t366 VDPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X48 VGND.t172 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 a_12310_25988# VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X49 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_12308_40142# a_12420_40104# VDPWR.t600 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X50 a_10108_28544.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 a_10958_27928.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X51 tdc_0.start_buffer_0.start_buff.t3 a_7140_10670# VGND.t263 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X52 VDPWR.t257 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t3 a_24240_17262# VDPWR.t256 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X53 VGND.t494 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t8 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t3 VGND.t493 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X54 a_25060_15196# variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VGND.t5 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X55 VGND.t244 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 a_12310_32834# VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X56 a_16292_6966# input_stage_0.fine_delay_unit_0.in a_16292_6702# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X57 VDPWR.t610 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t2 a_15680_14582# VDPWR.t609 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X58 a_10108_35390.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 a_10958_34774.t10 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X59 a_10108_30826.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X60 a_9330_15794# a_9330_15504# VDPWR.t193 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X61 VDPWR.t201 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VDPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X62 VDPWR.t239 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 VDPWR.t238 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X63 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t7 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t8 VGND.t507 VGND.t506 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X64 VGND.t226 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t4 a_25060_18144# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X65 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t4 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t9 VGND.t271 VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X66 VDPWR.t368 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t4 VDPWR.t367 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X67 a_10108_28544.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 a_10958_27928.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X68 a_24790_8050# input_stage_1.fine_delay_unit_1.in a_23820_8460# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X69 tdc_0.vernier_delay_line_0.stop_strong.t30 a_9330_16954.t10 VDPWR.t108 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X70 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t0 VDPWR.t621 VGND.t407 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X71 uo_out[0].t0 a_12310_23706# VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X72 a_10958_25646.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 a_10108_26262.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X73 a_24240_17262# variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t5 VDPWR.t259 VDPWR.t258 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X74 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 VDPWR.t104 VDPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X75 a_25060_26988# VGND.t344 variable_delay_short_0.variable_delay_unit_5.out VGND.t345 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X76 VDPWR.t91 tdc_0.start_buffer_0.start_buff.t11 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t6 VDPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X77 tdc_0.vernier_delay_line_0.stop_strong.t29 a_9330_16954.t11 VDPWR.t109 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X78 a_15680_14582# variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VDPWR.t612 VDPWR.t611 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X79 a_10958_34774.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 a_10108_35390.t4 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X80 uo_out[3].t1 a_12310_30552# VGND.t46 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X81 VGND.t245 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t2 a_16500_12516# VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X82 VGND.t78 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t8 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t2 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X83 VGND.t169 tdc_0.vernier_delay_line_0.stop_strong.t36 a_10958_32492.t11 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X84 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 VDPWR.t5 VDPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X85 VGND.t460 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t3 a_25060_26988# VGND.t459 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X86 VDPWR.t464 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t8 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t4 VDPWR.t463 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X87 VGND.t454 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t10 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t3 VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X88 a_10958_23364.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 a_10108_23452# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X89 VGND.t1 input_stage_0.fine_delay_unit_1.in a_16292_8344# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X90 VGND.t164 tdc_0.vernier_delay_line_0.stop_strong.t37 a_10958_39338.t6 VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X91 a_23820_7082# input_stage_1.fine_delay_unit_0.in a_24790_6672# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X92 VDPWR.t73 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t8 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t0 VDPWR.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X93 VDPWR.t190 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 VDPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X94 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X95 VGND.t165 tdc_0.vernier_delay_line_0.stop_strong.t38 a_10958_25646.t12 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X96 VGND.t496 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t6 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X97 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t1 ui_in[5].t1 VGND.t154 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X98 VDPWR.t561 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t7 VDPWR.t560 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X99 tdc_0.vernier_delay_line_0.stop_strong.t14 a_9330_16954.t12 VGND.t36 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X100 VDPWR.t396 tdc_0.vernier_delay_line_0.stop_strong.t39 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X101 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t9 VDPWR.t129 VDPWR.t128 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X102 a_10958_34774.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 a_10108_35390.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X103 a_13254_30598# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 uo_out[3].t2 VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X104 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t5 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t9 VDPWR.t220 VDPWR.t219 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X105 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t10 VGND.t300 VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X106 VGND.t335 tdc_0.vernier_delay_line_0.stop_strong.t40 a_10958_32492.t10 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X107 variable_delay_short_0.variable_delay_unit_5.forward.t1 variable_delay_short_0.variable_delay_unit_5.in.t2 VDPWR.t255 VDPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X108 a_9330_14344# a_9330_14054# VDPWR.t198 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X109 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 VGND.t341 VGND.t340 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X110 a_16292_8080# input_stage_0.fine_delay_unit_1.in a_15322_8490# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X111 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t3 tdc_0.start_buffer_0.start_buff.t12 VGND.t381 VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X112 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 a_10958_25646.t4 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X113 a_24790_6672# input_stage_1.fine_delay_unit_0.in a_23820_7082# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X114 a_9330_16954.t7 a_9330_15794# VDPWR.t599 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X115 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t7 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t8 VDPWR.t374 VDPWR.t373 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X116 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 VDPWR.t175 VDPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X117 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t0 VDPWR.t622 VGND.t406 VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X118 a_10958_23364.t4 tdc_0.vernier_delay_line_0.stop_strong.t41 VGND.t161 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X119 a_10108_30826.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 a_10958_30210.t8 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X120 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t0 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t9 VGND.t116 VGND.t115 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X121 a_25060_20210# ui_in[5].t2 VGND.t242 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X122 a_10958_30210.t4 tdc_0.vernier_delay_line_0.stop_strong.t42 VGND.t162 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X123 a_10108_23980.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 a_10958_23364.t10 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X124 variable_delay_short_0.variable_delay_unit_4.in.t1 variable_delay_short_0.variable_delay_unit_3.in.t2 VDPWR.t75 VDPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X125 VDPWR.t181 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t7 VDPWR.t180 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X126 a_15322_8490# input_stage_0.fine_delay_unit_1.in a_16292_8080# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X127 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t5 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t10 VGND.t505 VGND.t504 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X128 a_10958_39338.t5 tdc_0.vernier_delay_line_0.stop_strong.t43 VGND.t159 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X129 VDPWR.t297 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 VDPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X130 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t5 tdc_0.start_buffer_0.start_delay.t8 VDPWR.t36 VDPWR.t35 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X131 VDPWR.t275 ui_in[5].t3 a_24240_21092# VDPWR.t274 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X132 a_13254_24130# uo_out[0].t4 VGND.t110 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X133 VGND.t501 ui_in[5].t4 a_25060_20210# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X134 VGND.t309 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t4 VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X135 a_13254_33258# uo_out[4].t4 VGND.t532 VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X136 VGND.t160 tdc_0.vernier_delay_line_0.stop_strong.t44 a_10958_30210.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X137 a_16500_15464# variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t4 VGND.t59 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X138 a_24240_24040# ui_in[4].t0 VDPWR.t124 VDPWR.t123 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X139 VGND.t151 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X140 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 a_10958_34774.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X141 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 VDPWR.t113 VDPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X142 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 VDPWR.t541 VDPWR.t540 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X143 a_13254_40104# uo_out[7].t4 VGND.t241 VGND.t240 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X144 variable_delay_short_0.variable_delay_unit_5.forward.t0 variable_delay_short_0.variable_delay_unit_5.in.t3 VGND.t307 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X145 a_9330_15214# a_9330_14924# VGND.t203 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X146 a_24240_21092# ui_in[5].t5 VDPWR.t555 VDPWR.t554 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X147 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 VDPWR.t411 VDPWR.t410 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X148 VDPWR.t135 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12420_28316# VDPWR.t134 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X149 VGND.t189 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t0 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X150 a_25060_18144# variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.out VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X151 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t4 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t10 VGND.t175 VGND.t174 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X152 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 VDPWR.t127 VDPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X153 tdc_0.vernier_delay_line_0.stop_strong.t13 a_9330_16954.t13 VGND.t37 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X154 tdc_0.vernier_delay_line_0.start_pos.t7 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t8 VDPWR.t147 VDPWR.t146 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X155 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12308_37860# a_12420_37822# VDPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X156 VGND.t231 ui_in[7].t0 a_25060_14314# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X157 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 a_13254_30976# VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X158 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X159 tdc_0.vernier_delay_line_0.stop_strong.t12 a_9330_16954.t14 VGND.t38 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X160 VDPWR.t334 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 VDPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X161 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t6 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t10 VGND.t524 VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X162 a_24240_18144# ui_in[6].t0 VDPWR.t79 VDPWR.t78 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X163 tdc_0.vernier_delay_line_0.stop_strong.t11 a_9330_16954.t15 VGND.t35 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X164 a_25284_5108# ua[0].t0 VGND.t235 VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X165 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 VDPWR.t407 VDPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X166 VDPWR.t336 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VDPWR.t335 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X167 VGND.t202 uio_in[0].t0 a_25060_11366# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X168 variable_delay_short_0.variable_delay_unit_4.in.t0 variable_delay_short_0.variable_delay_unit_3.in.t3 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X169 VDPWR.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 VDPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X170 VGND.t465 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 VGND.t464 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X171 tdc_0.vernier_delay_line_0.stop_strong.t28 a_9330_16954.t16 VDPWR.t25 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X172 tdc_0.vernier_delay_line_0.start_neg.t5 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t8 VDPWR.t159 VDPWR.t158 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X173 a_24240_15196# ui_in[7].t1 VDPWR.t266 VDPWR.t265 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X174 VGND.t177 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t11 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t3 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X175 VDPWR.t97 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VDPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X176 VDPWR.t263 tdc_0.vernier_delay_line_0.start_pos.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 VDPWR.t262 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X177 VGND.t64 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_13254_39726# VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X178 a_15680_12516# VDPWR.t448 VDPWR.t450 VDPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X179 VGND.t370 tdc_0.start_buffer_0.start_delay.t9 tdc_0.start_buffer_0.start_buff.t9 VGND.t369 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X180 VDPWR.t163 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 VDPWR.t162 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X181 a_10108_33108.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 a_10958_32492.t4 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X182 VDPWR.t81 ui_in[6].t1 a_24240_18144# VDPWR.t80 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X183 a_25060_26106# VDPWR.t623 VGND.t405 VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X184 VDPWR.t251 tdc_0.start_buffer_0.start_buff.t13 tdc_0.start_buffer_0.start_delay.t5 VDPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X185 variable_delay_dummy_0.variable_delay_unit_1.forward.t0 variable_delay_dummy_0.variable_delay_unit_1.in.t2 VGND.t305 VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X186 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X187 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 VDPWR.t402 VDPWR.t401 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X188 a_9330_13764# variable_delay_short_0.out VGND.t544 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X189 VDPWR.t447 VDPWR.t445 a_15680_15464# VDPWR.t446 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X190 VGND.t339 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 VGND.t338 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X191 VGND.t53 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X192 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 VDPWR.t490 VDPWR.t489 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X193 a_24240_26988# VGND.t562 variable_delay_short_0.variable_delay_unit_5.out VDPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X194 VDPWR.t188 tdc_0.vernier_delay_line_0.stop_strong.t45 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VDPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X195 a_25060_23158# ui_in[4].t1 VGND.t108 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X196 VDPWR.t142 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t7 VDPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X197 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VDPWR.t192 VDPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X198 VGND.t353 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X199 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 VDPWR.t391 VDPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X200 VDPWR.t444 VDPWR.t442 a_24240_26988# VDPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X201 VDPWR.t34 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t9 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t1 VDPWR.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X202 a_10958_30210.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 a_10108_30826.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X203 tdc_0.start_buffer_0.start_buff.t7 a_7140_10670# VDPWR.t304 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X204 a_23820_7082# input_stage_1.fine_delay_unit_0.in VDPWR.t462 VDPWR.t461 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X205 a_16786_5138# ua[0].t1 VGND.t237 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X206 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 VDPWR.t333 VDPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X207 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.start_pos.t9 VGND.t66 VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X208 VDPWR.t618 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12420_37444# VDPWR.t617 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X209 a_24790_8314# ui_in[2].t0 a_24790_8050# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X210 VDPWR.t518 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t1 VDPWR.t517 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X211 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 VGND.t55 VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X212 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 VGND.t448 VGND.t447 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X213 tdc_0.start_buffer_0.start_buff.t2 a_7140_10670# VGND.t262 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X214 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 VGND.t357 VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X215 VDPWR.t499 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 VDPWR.t498 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X216 VDPWR.t99 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X217 tdc_0.start_buffer_0.start_delay.t7 tdc_0.start_buffer_0.start_buff.t14 VGND.t379 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X218 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 VDPWR.t393 VDPWR.t392 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X219 a_12420_26412# uo_out[1].t4 VDPWR.t295 VDPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X220 a_9330_15214# a_9330_14924# VDPWR.t225 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X221 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t4 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t10 VGND.t122 VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X222 VGND.t327 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X223 tdc_0.vernier_delay_line_0.start_pos.t4 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t10 VGND.t528 VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X224 VGND.t456 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X225 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.start_neg.t8 VDPWR.t161 VDPWR.t160 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X226 a_24240_20210# variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t4 VDPWR.t354 VDPWR.t353 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X227 tdc_0.vernier_delay_line_0.stop_strong.t27 a_9330_16954.t17 VDPWR.t26 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X228 VDPWR.t481 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 VDPWR.t480 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X229 a_15322_8490# input_stage_0.fine_delay_unit_1.in VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X230 VGND.t291 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t2 VGND.t290 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X231 VGND.t158 tdc_0.vernier_delay_line_0.stop_strong.t46 a_10958_37056.t9 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X232 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 a_10958_30210.t12 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X233 tdc_0.vernier_delay_line_0.stop_strong.t26 a_9330_16954.t18 VDPWR.t23 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X234 tdc_0.vernier_delay_line_0.start_neg.t2 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t10 VGND.t140 VGND.t139 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X235 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 VDPWR.t329 VDPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X236 VDPWR.t338 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 a_12310_28270# VDPWR.t337 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X237 variable_delay_dummy_0.in a_15322_8490# VDPWR.t166 VDPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X238 VGND.t403 VDPWR.t624 a_16500_14582# VGND.t402 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X239 tdc_0.vernier_delay_line_0.stop_strong.t25 a_9330_16954.t19 VDPWR.t24 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X240 a_12420_32880# a_12310_32834# uo_out[4].t1 VDPWR.t194 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X241 VGND.t157 tdc_0.vernier_delay_line_0.stop_strong.t47 a_10958_27928.t8 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X242 VGND.t80 tdc_0.vernier_delay_line_0.start_pos.t10 tdc_0.vernier_delay_line_0.start_neg.t6 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X243 VDPWR.t38 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 a_12310_37398# VDPWR.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X244 a_13254_28316# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 uo_out[2].t0 VGND.t349 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X245 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t48 VDPWR.t186 VDPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X246 a_16292_8344# uio_in[3].t0 a_16292_8080# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X247 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 VGND.t389 VGND.t388 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X248 a_24790_6936# ui_in[0].t0 a_24790_6672# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X249 VDPWR.t356 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t5 a_24240_20210# VDPWR.t355 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X250 a_13254_37822# uo_out[6].t4 VGND.t321 VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X251 input_stage_0.fine_delay_unit_0.in input_stage_0.nand_gate_0.out VDPWR.t608 VDPWR.t607 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X252 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.stop_strong.t49 VDPWR.t381 VDPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X253 VDPWR.t614 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12420_23752# VDPWR.t613 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X254 a_16500_14582# VDPWR.t625 VGND.t401 VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X255 VDPWR.t567 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12420_32880# VDPWR.t566 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X256 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 a_13254_28694# VGND.t238 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X257 a_10958_25646.t11 tdc_0.vernier_delay_line_0.stop_strong.t50 VGND.t317 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X258 VGND.t561 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 a_12310_39680# VGND.t560 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X259 VDPWR.t117 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VDPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X260 a_9330_13764# variable_delay_short_0.out VDPWR.t605 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X261 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 a_10108_39426# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X262 uo_out[5].t0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t347 VDPWR.t346 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X263 VGND.t477 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_13254_26034# VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X264 VDPWR.t119 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X265 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t0 ui_in[6].t2 VDPWR.t306 VDPWR.t305 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X266 a_10108_37672.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X267 a_24240_18144# variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.out VDPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X268 VDPWR.t276 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 VDPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X269 VDPWR.t406 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t4 a_24240_14314# VDPWR.t405 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X270 a_15680_15464# VGND.t563 variable_delay_dummy_0.variable_delay_unit_1.out VDPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X271 a_25060_12248# variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t3 VGND.t292 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X272 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t0 ui_in[7].t2 VDPWR.t533 VDPWR.t527 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X273 a_12420_26034# a_12310_25988# uo_out[1].t0 VDPWR.t195 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X274 VGND.t57 tdc_0.vernier_delay_line_0.start_neg.t9 tdc_0.vernier_delay_line_0.start_pos.t0 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X275 VDPWR.t278 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t3 a_15680_11634# VDPWR.t277 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X276 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 a_10108_28544.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X277 uo_out[7].t3 a_12310_39680# VGND.t85 VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X278 a_12420_35540# uo_out[5].t4 VDPWR.t483 VDPWR.t482 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X279 VDPWR.t342 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t4 a_24240_11366# VDPWR.t341 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X280 VDPWR.t466 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VDPWR.t465 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X281 VGND.t387 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 VGND.t386 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X282 VGND.t83 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X283 VDPWR.t458 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 VDPWR.t457 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X284 a_10108_28016# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X285 VGND.t517 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t11 tdc_0.vernier_delay_line_0.start_pos.t3 VGND.t516 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X286 VDPWR.t395 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 a_12310_23706# VDPWR.t394 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X287 a_10958_39338.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 a_10108_39426# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X288 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.start_neg.t10 VGND.t303 VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X289 a_24240_26106# variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t4 VDPWR.t509 VDPWR.t508 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X290 VGND.t153 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X291 VDPWR.t69 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 a_12310_30552# VDPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X292 tdc_0.vernier_delay_line_0.stop_strong.t10 a_9330_16954.t20 VGND.t34 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X293 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 VGND.t285 VGND.t284 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X294 VDPWR.t314 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t11 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t2 VDPWR.t313 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X295 VGND.t359 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t4 a_25060_24040# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X296 a_13254_37444# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 uo_out[6].t1 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X297 a_24240_23158# variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t5 VDPWR.t203 VDPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X298 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VGND.t225 VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X299 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t6 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t11 VDPWR.t559 VDPWR.t558 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X300 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 a_10108_25734# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X301 VGND.t223 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t6 a_25060_21092# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X302 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 VGND.t147 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X303 a_10108_23980.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X304 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t1 ui_in[6].t3 VGND.t264 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X305 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t7 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t11 VDPWR.t497 VDPWR.t496 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X306 a_10958_39338.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 a_10108_39426# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X307 a_10108_37672.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 a_10958_37056.t11 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X308 VGND.t206 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 a_12310_35116# VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X309 variable_delay_short_0.variable_delay_unit_5.in.t0 variable_delay_short_0.variable_delay_unit_4.in.t2 VDPWR.t71 VDPWR.t70 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X310 a_10958_34774.t8 tdc_0.vernier_delay_line_0.stop_strong.t51 VGND.t217 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X311 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 VGND.t413 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X312 VDPWR.t563 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VDPWR.t562 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X313 input_stage_0.fine_delay_unit_1.in a_15322_7112# VDPWR.t415 VDPWR.t414 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X314 VGND.t325 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13254_35162# VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X315 input_stage_1.fine_delay_unit_1.in a_23820_7082# VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X316 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t1 ui_in[7].t3 VGND.t482 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X317 tdc_0.vernier_delay_line_0.stop_strong.t9 a_9330_16954.t21 VGND.t32 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X318 VDPWR.t616 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t10 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t4 VDPWR.t615 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X319 a_10958_27928.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 a_10108_28544.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X320 uo_out[1].t1 a_12310_25988# VGND.t182 VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X321 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t0 VDPWR.t626 VGND.t399 VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X322 VDPWR.t213 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VDPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X323 tdc_0.vernier_delay_line_0.stop_strong.t8 a_9330_16954.t22 VGND.t33 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X324 VDPWR.t310 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t6 VDPWR.t309 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X325 a_10108_37672.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 a_10958_37056.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X326 a_12420_30976# uo_out[3].t4 VDPWR.t211 VDPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X327 input_stage_1.nand_gate_0.out ua[0].t2 VDPWR.t534 VDPWR.t426 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X328 VGND.t4 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t5 a_25060_15196# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X329 uo_out[4].t2 a_12310_32834# VGND.t180 VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X330 VGND.t411 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X331 VDPWR.t144 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t10 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t7 VDPWR.t143 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X332 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 a_10108_30826.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X333 a_10108_28016# tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 a_10958_27928.t12 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X334 variable_delay_short_0.variable_delay_unit_3.in.t1 variable_delay_short_0.variable_delay_unit_2.in.t2 VDPWR.t549 VDPWR.t305 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X335 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 VDPWR.t155 VDPWR.t154 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X336 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t3 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t11 VDPWR.t364 VDPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X337 a_10958_27928.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 a_10108_28544.t4 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X338 a_24790_8314# input_stage_1.fine_delay_unit_1.in a_24790_8050# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X339 a_13254_23752# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 uo_out[0].t2 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X340 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 VDPWR.t106 VDPWR.t105 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X341 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 VDPWR.t399 VDPWR.t398 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X342 VGND.t429 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t6 VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X343 a_10958_32492.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 a_10108_32580# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X344 variable_delay_short_0.variable_delay_unit_2.in.t0 variable_delay_short_0.variable_delay_unit_1.in.t2 VDPWR.t528 VDPWR.t527 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X345 a_10958_37056.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 a_10108_37672.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X346 a_16292_6702# input_stage_0.fine_delay_unit_0.in a_15322_7112# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X347 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t5 tdc_0.start_buffer_0.start_buff.t15 VDPWR.t253 VDPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X348 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.forward.t2 a_15680_14582# VDPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X349 a_9330_14634# a_9330_14344# VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X350 VGND.t218 tdc_0.vernier_delay_line_0.stop_strong.t52 a_10958_34774.t7 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X351 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t1 VDPWR.t440 VDPWR.t441 VDPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X352 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t1 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t11 VGND.t253 VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X353 a_16500_12516# variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t4 VGND.t497 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X354 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 a_13254_24130# VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X355 a_10958_25646.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 a_10108_25734# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X356 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t5 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t11 VDPWR.t488 VDPWR.t487 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X357 a_10108_23980.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 a_10958_23364.t8 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X358 a_9330_16954.t2 a_9330_15794# VGND.t539 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X359 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t13 VGND.t269 VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X360 a_10108_33108.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X361 tdc_0.start_buffer_0.start_buff.t6 a_7140_10670# VDPWR.t303 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X362 a_10108_28016# tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 a_10958_27928.t11 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X363 VGND.t61 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t5 a_16500_15464# VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X364 variable_delay_short_0.variable_delay_unit_5.in.t1 variable_delay_short_0.variable_delay_unit_4.in.t3 VGND.t138 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X365 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 a_10108_34862# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X366 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t11 VGND.t124 VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X367 tdc_0.start_buffer_0.start_delay.t4 tdc_0.start_buffer_0.start_buff.t16 VDPWR.t172 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X368 a_25060_15196# variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_1.out VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X369 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t0 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t12 VDPWR.t261 VDPWR.t260 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X370 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 a_10958_34774.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X371 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 a_10108_23980.t4 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X372 input_stage_0.nand_gate_0.out ua[0].t3 VDPWR.t535 VDPWR.t531 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X373 a_10958_32492.t9 tdc_0.vernier_delay_line_0.stop_strong.t53 VGND.t91 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X374 VGND.t216 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_13254_30598# VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X375 tdc_0.vernier_delay_line_0.stop_strong.t24 a_9330_16954.t23 VDPWR.t22 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X376 VGND.t432 input_stage_0.fine_delay_unit_0.in a_16292_6966# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X377 a_25060_12248# variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.out VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X378 tdc_0.start_buffer_0.start_buff.t1 a_7140_10670# VGND.t261 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X379 VGND.t208 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X380 VDPWR.t140 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t6 VDPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X381 a_10958_25646.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 a_10108_25734# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X382 a_24790_6936# input_stage_1.fine_delay_unit_0.in a_24790_6672# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X383 VGND.t323 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t5 VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X384 VDPWR.t177 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 VDPWR.t176 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X385 VGND.t92 tdc_0.vernier_delay_line_0.stop_strong.t54 a_10958_23364.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X386 variable_delay_short_0.variable_delay_unit_3.in.t0 variable_delay_short_0.variable_delay_unit_2.in.t3 VGND.t265 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X387 a_25060_24040# variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_4.out VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X388 VGND.t313 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 VGND.t312 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X389 a_10958_30210.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 a_10108_30826.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X390 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X391 a_24240_12248# uio_in[0].t1 VDPWR.t222 VDPWR.t221 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X392 a_12420_39726# a_12310_39680# uo_out[7].t2 VDPWR.t85 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X393 VGND.t462 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t5 a_25060_26988# VGND.t461 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X394 VDPWR.t209 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t12 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t1 VDPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X395 variable_delay_short_0.variable_delay_unit_2.in.t1 variable_delay_short_0.variable_delay_unit_1.in.t3 VGND.t475 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X396 a_10958_23364.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 a_10108_23980.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X397 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t6 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t12 VDPWR.t468 VDPWR.t467 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X398 tdc_0.vernier_delay_line_0.stop_strong.t23 a_9330_16954.t24 VDPWR.t20 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X399 a_16292_8080# input_stage_0.fine_delay_unit_1.in a_15322_8490# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X400 VGND.t99 tdc_0.vernier_delay_line_0.stop_strong.t55 a_10958_39338.t4 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X401 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 VGND.t210 VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X402 variable_delay_dummy_0.variable_delay_unit_1.in.t0 variable_delay_dummy_0.in VGND.t512 VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X403 tdc_0.vernier_delay_line_0.stop_strong.t22 a_9330_16954.t25 VDPWR.t21 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X404 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.stop_strong.t56 VDPWR.t114 VDPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X405 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 VDPWR.t288 VDPWR.t287 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X406 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X407 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t5 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t11 VDPWR.t501 VDPWR.t500 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X408 a_25060_20210# ui_in[5].t6 VGND.t500 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X409 a_10108_33108.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 a_10958_32492.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X410 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 a_13254_33258# VGND.t508 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X411 a_10958_30210.t2 tdc_0.vernier_delay_line_0.stop_strong.t57 VGND.t195 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X412 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t11 VGND.t118 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X413 VDPWR.t121 ui_in[4].t2 a_24240_24040# VDPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X414 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 VGND.t334 VGND.t333 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X415 a_10958_34774.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 a_10108_34862# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X416 VDPWR.t492 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 VDPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X417 VDPWR.t470 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t13 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t5 VDPWR.t469 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X418 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t2 tdc_0.start_buffer_0.start_buff.t17 VGND.t378 VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X419 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t170 VDPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X420 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 a_13254_40104# VGND.t193 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X421 a_10958_23364.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 a_10108_23980.t0 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X422 VDPWR.t404 tdc_0.start_buffer_0.start_delay.t10 tdc_0.start_buffer_0.start_buff.t8 VDPWR.t403 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X423 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t13 VGND.t331 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X424 VDPWR.t553 ui_in[5].t7 a_24240_21092# VDPWR.t552 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X425 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t348 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X426 VGND.t287 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t6 a_25060_18144# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X427 variable_delay_dummy_0.variable_delay_unit_1.forward.t1 variable_delay_dummy_0.variable_delay_unit_1.in.t3 VDPWR.t138 VDPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X428 a_9330_14634# a_9330_14344# VDPWR.t164 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X429 a_24790_8050# input_stage_1.fine_delay_unit_1.in a_23820_8460# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X430 a_25060_14314# ui_in[7].t4 VGND.t518 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X431 VDPWR.t31 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 VDPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X432 VGND.t149 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X433 VDPWR.t370 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 VDPWR.t369 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X434 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X435 VGND.t48 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t12 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t0 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X436 a_9330_16954.t6 a_9330_15794# VDPWR.t598 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X437 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 a_10108_39954.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X438 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 a_10958_37056.t4 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X439 input_stage_1.nand_gate_0.out VDPWR.t627 a_25284_5108# VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X440 VDPWR.t216 tdc_0.vernier_delay_line_0.stop_strong.t58 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 VDPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X441 VGND.t214 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t12 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t0 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X442 a_25060_11366# uio_in[0].t2 VGND.t131 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X443 variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_3.in.t4 a_25060_17262# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X444 VDPWR.t207 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 VDPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X445 VGND.t228 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t13 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t1 VGND.t227 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X446 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 VGND.t441 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X447 VDPWR.t286 tdc_0.vernier_delay_line_0.stop_strong.t59 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X448 VDPWR.t576 ui_in[7].t5 a_24240_15196# VDPWR.t575 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X449 a_23820_8460# input_stage_1.fine_delay_unit_1.in a_24790_8050# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X450 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.in.t4 a_25060_14314# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X451 a_16500_15464# VGND.t342 variable_delay_dummy_0.variable_delay_unit_1.out VGND.t343 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X452 VGND.t279 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t12 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t2 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X453 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 tdc_0.vernier_delay_line_0.start_pos.t11 VDPWR.t299 VDPWR.t298 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X454 VDPWR.t439 VDPWR.t437 a_15680_12516# VDPWR.t438 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X455 a_10958_32492.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 a_10108_33108.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X456 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 VDPWR.t372 VDPWR.t371 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X457 VGND.t398 VDPWR.t628 a_16500_11634# VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X458 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t2 tdc_0.start_buffer_0.start_delay.t11 VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X459 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 VDPWR.t183 VDPWR.t182 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X460 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.forward.t2 a_25060_26106# VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X461 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 VDPWR.t93 VDPWR.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X462 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 a_10108_30298# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X463 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 VGND.t44 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X464 uo_out[2].t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t537 VDPWR.t536 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X465 tdc_0.vernier_delay_line_0.stop_strong.t7 a_9330_16954.t26 VGND.t31 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X466 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t6 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t12 VDPWR.t316 VDPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X467 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 VGND.t247 VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X468 VDPWR.t60 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 VDPWR.t59 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X469 VGND.t366 tdc_0.start_buffer_0.start_delay.t12 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t1 VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X470 a_10108_30298# tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 a_10958_30210.t11 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X471 VDPWR.t505 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 VDPWR.t504 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X472 tdc_0.vernier_delay_line_0.start_pos.t6 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t12 VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X473 a_10108_35390.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 a_10958_34774.t12 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X474 VDPWR.t269 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t4 VDPWR.t268 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X475 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t157 VDPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X476 a_12420_28694# uo_out[2].t4 VDPWR.t325 VDPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X477 VGND.t362 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X478 VGND.t479 ui_in[3].t0 a_24790_8314# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X479 tdc_0.vernier_delay_line_0.start_neg.t4 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t11 VDPWR.t376 VDPWR.t375 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X480 VGND.t355 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 VGND.t354 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X481 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 a_10958_23364.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X482 a_24240_15196# variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_1.out VDPWR.t61 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X483 VGND.t76 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X484 a_10958_39338.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 a_10108_39954.t3 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X485 VDPWR.t50 tdc_0.vernier_delay_line_0.start_pos.t12 tdc_0.vernier_delay_line_0.start_neg.t7 VDPWR.t49 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X486 a_15680_12516# variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.out VDPWR.t548 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X487 a_16292_6966# uio_in[1].t0 a_16292_6702# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X488 VGND.t135 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X489 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 VDPWR.t87 VDPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X490 a_10958_30210.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 a_10108_30298# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X491 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t0 uio_in[0].t3 VDPWR.t151 VDPWR.t150 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X492 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 VDPWR.t235 VDPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X493 a_25060_26106# VDPWR.t629 VGND.t397 VGND.t396 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X494 a_24240_12248# variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.out VDPWR.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X495 VGND.t120 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X496 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12308_26450# a_12420_26412# VDPWR.t264 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X497 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t0 ui_in[4].t3 VDPWR.t122 VDPWR.t70 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X498 a_24240_24040# variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_4.out VDPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X499 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 VGND.t70 VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X500 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 VGND.t557 VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X501 a_25060_23158# ui_in[4].t4 VGND.t525 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X502 VGND.t254 tdc_0.vernier_delay_line_0.stop_strong.t60 a_10958_37056.t8 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X503 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t61 VDPWR.t215 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X504 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12308_35578# a_12420_35540# VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X505 VDPWR.t436 VDPWR.t434 a_24240_26988# VDPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X506 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 VGND.t418 VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X507 a_10958_30210.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 a_10108_30298# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X508 VGND.t201 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t12 tdc_0.vernier_delay_line_0.start_neg.t1 VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X509 a_9330_14054# a_9330_13764# VGND.t515 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X510 a_10958_27928.t7 tdc_0.vernier_delay_line_0.stop_strong.t62 VGND.t194 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X511 VDPWR.t345 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VDPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X512 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 tdc_0.vernier_delay_line_0.start_pos.t13 VGND.t436 VGND.t435 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X513 uo_out[6].t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t620 VDPWR.t619 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X514 VGND.t112 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_13254_28316# VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X515 input_stage_1.fine_delay_unit_0.in input_stage_1.nand_gate_0.out VGND.t133 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X516 a_9330_15504# a_9330_15214# VGND.t348 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X517 a_10108_39954.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X518 VGND.t480 uio_in[4].t0 a_16292_8344# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X519 VDPWR.t133 tdc_0.vernier_delay_line_0.start_neg.t11 tdc_0.vernier_delay_line_0.start_pos.t1 VDPWR.t132 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X520 a_9330_16954.t1 a_9330_15794# VGND.t538 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X521 a_24240_20210# variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t7 VDPWR.t245 VDPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X522 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 a_13254_37822# VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X523 a_25060_17262# ui_in[6].t4 VGND.t62 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X524 tdc_0.vernier_delay_line_0.stop_strong.t6 a_9330_16954.t27 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X525 VDPWR.t168 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 VDPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X526 tdc_0.start_buffer_0.start_buff.t5 a_7140_10670# VDPWR.t302 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X527 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.forward.t3 a_16500_14582# VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X528 VGND.t212 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X529 tdc_0.vernier_delay_line_0.stop_strong.t5 a_9330_16954.t28 VGND.t30 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X530 VDPWR.t11 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t13 tdc_0.vernier_delay_line_0.start_pos.t5 VDPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X531 VGND.t233 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X532 VGND.t468 tdc_0.vernier_delay_line_0.stop_strong.t63 a_10958_25646.t10 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X533 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t3 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t13 VGND.t534 VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X534 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t41 VDPWR.t40 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X535 a_12420_35162# a_12310_35116# uo_out[5].t3 VDPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X536 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t1 uio_in[0].t4 VGND.t439 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X537 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 a_10108_37672.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X538 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.start_neg.t12 VDPWR.t224 VDPWR.t223 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X539 VGND.t469 tdc_0.vernier_delay_line_0.stop_strong.t64 a_10958_34774.t6 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X540 tdc_0.start_buffer_0.start_buff.t0 a_7140_10670# VGND.t260 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X541 VDPWR.t52 ui_in[6].t5 a_24240_18144# VDPWR.t51 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X542 tdc_0.vernier_delay_line_0.stop_strong.t21 a_9330_16954.t29 VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X543 VGND.t337 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VGND.t336 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X544 VDPWR.t280 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 VDPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X545 VDPWR.t573 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 a_12310_25988# VDPWR.t572 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X546 a_24240_14314# variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VDPWR.t95 VDPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X547 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t1 ui_in[4].t5 VGND.t526 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X548 VGND.t420 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X549 tdc_0.start_buffer_0.start_delay.t2 tdc_0.start_buffer_0.start_buff.t18 VGND.t376 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X550 VDPWR.t433 VDPWR.t431 a_15680_15464# VDPWR.t432 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X551 VGND.t535 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t5 a_25060_12248# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X552 a_15680_11634# variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t5 VDPWR.t547 VDPWR.t546 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X553 VDPWR.t565 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 a_12310_32834# VDPWR.t564 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X554 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 VGND.t484 VGND.t483 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X555 variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_3.in.t5 a_24240_17262# VDPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X556 a_24240_11366# variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t6 VDPWR.t593 VDPWR.t592 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X557 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 VDPWR.t507 VDPWR.t506 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X558 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 VGND.t385 VGND.t384 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X559 a_23820_8460# input_stage_1.fine_delay_unit_1.in VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X560 VGND.t458 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 VGND.t457 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X561 variable_delay_short_0.in a_23820_8460# VDPWR.t77 VDPWR.t76 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X562 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 VGND.t514 VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X563 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 VDPWR.t456 VDPWR.t455 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X564 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.in.t5 a_24240_14314# VDPWR.t516 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X565 uo_out[0].t3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t318 VDPWR.t317 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X566 variable_delay_short_0.variable_delay_unit_1.in.t1 variable_delay_short_0.in VDPWR.t300 VDPWR.t150 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X567 VGND.t68 tdc_0.vernier_delay_line_0.start_neg.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X568 variable_delay_dummy_0.out variable_delay_dummy_0.variable_delay_unit_1.in.t4 a_15680_11634# VDPWR.t115 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X569 a_10108_39954.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 a_10958_39338.t9 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X570 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.forward.t3 a_24240_26106# VDPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X571 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t1 VDPWR.t428 VDPWR.t430 VDPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X572 variable_delay_dummy_0.in a_15322_8490# VGND.t143 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X573 uo_out[3].t3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t539 VDPWR.t538 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X574 a_10958_25646.t9 tdc_0.vernier_delay_line_0.stop_strong.t65 VGND.t452 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X575 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 VGND.t249 VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X576 input_stage_1.fine_delay_unit_0.in input_stage_1.nand_gate_0.out VDPWR.t153 VDPWR.t152 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X577 VGND.t555 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_13254_37444# VGND.t554 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X578 VGND.t315 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 VGND.t314 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X579 VDPWR.t454 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 VDPWR.t453 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X580 a_10108_39954.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 a_10958_39338.t8 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X581 a_10958_37056.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 a_10108_37672.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X582 a_12420_30598# a_12310_30552# uo_out[3].t0 VDPWR.t32 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X583 a_9330_14054# a_9330_13764# VDPWR.t574 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X584 a_13254_26412# uo_out[1].t5 VGND.t257 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X585 VDPWR.t472 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t13 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t7 VDPWR.t471 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X586 VGND.t137 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X587 a_9330_15504# a_9330_15214# VDPWR.t400 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X588 a_9330_16954.t5 a_9330_15794# VDPWR.t597 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X589 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t3 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t13 VDPWR.t495 VDPWR.t494 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X590 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.stop_strong.t66 VDPWR.t493 VDPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X591 tdc_0.vernier_delay_line_0.stop_strong.t20 a_9330_16954.t30 VDPWR.t110 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X592 a_25060_21092# variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.out VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X593 VGND.t486 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 a_12310_28270# VGND.t485 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X594 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t5 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t14 VDPWR.t308 VDPWR.t307 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X595 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 a_10108_28016# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X596 a_24240_26106# variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t6 VDPWR.t243 VDPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X597 VGND.t470 tdc_0.vernier_delay_line_0.stop_strong.t67 a_10958_37056.t7 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X598 a_13254_32880# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 uo_out[4].t3 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X599 a_10108_26262.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X600 VDPWR.t427 VDPWR.t425 input_stage_1.nand_gate_0.out VDPWR.t426 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X601 tdc_0.vernier_delay_line_0.stop_strong.t19 a_9330_16954.t31 VDPWR.t111 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X602 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t6 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t13 VDPWR.t387 VDPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X603 VGND.t190 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t6 a_25060_24040# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X604 VGND.t74 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 a_12310_37398# VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X605 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 VGND.t409 VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X606 variable_delay_short_0.variable_delay_unit_1.in.t0 variable_delay_short_0.in VGND.t258 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X607 a_24240_23158# variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t7 VDPWR.t205 VDPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X608 VGND.t27 input_stage_1.fine_delay_unit_1.in a_24790_8314# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X609 VGND.t549 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_13254_23752# VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X610 a_12420_24130# uo_out[0].t5 VDPWR.t131 VDPWR.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X611 VDPWR.t65 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 VDPWR.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X612 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 a_10958_37056.t5 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X613 a_15322_7112# input_stage_0.fine_delay_unit_0.in a_16292_6702# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X614 VGND.t510 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_13254_32880# VGND.t509 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X615 tdc_0.vernier_delay_line_0.stop_strong.t4 a_9330_16954.t32 VGND.t97 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X616 a_10958_34774.t5 tdc_0.vernier_delay_line_0.stop_strong.t68 VGND.t471 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X617 VGND.t316 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t6 a_16500_12516# VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X618 VDPWR.t323 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t14 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t3 VDPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X619 a_12420_33258# uo_out[4].t5 VDPWR.t589 VDPWR.t588 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X620 VDPWR.t360 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 VDPWR.t359 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X621 VGND.t184 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X622 uo_out[5].t2 a_12310_35116# VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X623 a_10108_26262.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 a_10958_25646.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X624 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 a_10108_33108.t5 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X625 a_10958_27928.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 a_10108_28016# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X626 a_12420_40104# uo_out[7].t5 VDPWR.t273 VDPWR.t272 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X627 a_24240_17262# variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t7 VDPWR.t327 VDPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X628 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 VDPWR.t67 VDPWR.t66 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X629 a_13254_26034# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 uo_out[1].t2 VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X630 a_16292_6702# input_stage_0.fine_delay_unit_0.in a_15322_7112# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X631 a_15680_14582# variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VDPWR.t485 VDPWR.t484 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X632 VGND.t3 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t7 a_25060_15196# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X633 a_10958_34774.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 a_10108_34862# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X634 variable_delay_dummy_0.variable_delay_unit_1.in.t1 variable_delay_dummy_0.in VDPWR.t569 VDPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X635 a_13254_35540# uo_out[5].t5 VGND.t126 VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X636 VGND.t93 tdc_0.vernier_delay_line_0.stop_strong.t69 a_10958_32492.t8 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X637 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12308_31014# a_12420_30976# VDPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X638 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 VDPWR.t13 VDPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X639 a_10958_25646.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 a_10108_26262.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X640 input_stage_0.fine_delay_unit_1.in a_15322_7112# VGND.t360 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X641 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t14 VGND.t422 VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X642 VGND.t267 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t0 VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X643 VGND.t536 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t7 a_25060_12248# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X644 a_15680_11634# variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t7 VDPWR.t380 VDPWR.t379 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X645 a_10958_27928.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 a_10108_28016# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X646 a_10108_26262.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 a_10958_25646.t0 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X647 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t5 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t13 VDPWR.t321 VDPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X648 VGND.t329 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 a_12310_23706# VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X649 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 VDPWR.t551 VDPWR.t550 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X650 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t4 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t15 VGND.t281 VGND.t280 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X651 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 VGND.t298 VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X652 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 a_10108_37144# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X653 VGND.t94 tdc_0.vernier_delay_line_0.stop_strong.t70 a_10958_30210.t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X654 VDPWR.t478 uio_in[0].t5 a_24240_12248# VDPWR.t477 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X655 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t4 tdc_0.start_buffer_0.start_buff.t19 VDPWR.t249 VDPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X656 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t1 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t14 VGND.t444 VGND.t443 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X657 VGND.t551 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 a_12310_30552# VGND.t550 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X658 a_16500_12516# variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.out VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X659 a_10958_32492.t7 tdc_0.vernier_delay_line_0.stop_strong.t71 VGND.t425 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X660 VDPWR.t58 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_12420_39726# VDPWR.t57 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X661 a_25060_26988# variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t7 VGND.t222 VGND.t221 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X662 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t2 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t14 VDPWR.t237 VDPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X663 a_10108_23452# tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 a_10958_23364.t12 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X664 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_5.in.t4 a_25060_23158# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X665 a_16292_8344# input_stage_0.fine_delay_unit_1.in a_16292_8080# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X666 a_10958_39338.t3 tdc_0.vernier_delay_line_0.stop_strong.t72 VGND.t427 VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X667 a_24790_6672# input_stage_1.fine_delay_unit_0.in a_23820_7082# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X668 VDPWR.t580 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 VDPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X669 a_9330_14924# a_9330_14634# VGND.t255 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X670 VGND.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X671 VDPWR.t271 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t13 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t4 VDPWR.t270 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X672 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t293 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X673 input_stage_0.nand_gate_0.out uio_in[5].t0 a_16786_5138# VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X674 VGND.t446 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t0 VGND.t445 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X675 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_4.in.t4 a_25060_20210# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X676 a_10958_32492.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 a_10108_33108.t0 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X677 VDPWR.t520 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t14 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t1 VDPWR.t519 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X678 VGND.t434 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X679 VGND.t442 tdc_0.vernier_delay_line_0.stop_strong.t73 a_10958_30210.t0 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X680 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X681 a_9330_16954.t0 a_9330_15794# VGND.t537 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X682 VDPWR.t557 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t14 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t4 VDPWR.t556 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X683 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 VDPWR.t232 VDPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X684 tdc_0.start_buffer_0.start_buff.t4 a_7140_10670# VDPWR.t301 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X685 VDPWR.t479 tdc_0.vernier_delay_line_0.stop_strong.t74 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X686 VGND.t375 tdc_0.start_buffer_0.start_buff.t20 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t1 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X687 VDPWR.t543 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t14 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t3 VDPWR.t542 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X688 tdc_0.vernier_delay_line_0.stop_strong.t3 a_9330_16954.t33 VGND.t39 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X689 tdc_0.start_buffer_0.start_delay.t3 tdc_0.start_buffer_0.start_buff.t21 VDPWR.t284 VDPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X690 tdc_0.vernier_delay_line_0.stop_strong.t2 a_9330_16954.t34 VGND.t40 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X691 VGND.t543 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X692 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X693 VGND.t251 tdc_0.vernier_delay_line_0.stop_strong.t75 a_10958_23364.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X694 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t4 tdc_0.start_buffer_0.start_delay.t13 VDPWR.t46 VDPWR.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X695 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 VGND.t18 VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X696 VGND.t199 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t1 VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X697 a_13254_30976# uo_out[3].t5 VGND.t192 VGND.t191 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X698 tdc_0.vernier_delay_line_0.stop_strong.t18 a_9330_16954.t35 VDPWR.t27 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X699 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 tdc_0.vernier_delay_line_0.stop_strong.t76 VDPWR.t285 VDPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X700 VGND.t431 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t14 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t7 VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X701 VGND.t499 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 VGND.t498 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X702 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 VDPWR.t522 VDPWR.t521 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X703 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 VGND.t488 VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X704 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 a_10108_23452# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X705 tdc_0.start_buffer_0.start_delay.t1 tdc_0.start_buffer_0.start_buff.t22 VGND.t373 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X706 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t7 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t15 VGND.t559 VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X707 VGND.t503 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t6 VGND.t502 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X708 a_10958_37056.t12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 a_10108_37144# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X709 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 VGND.t473 VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X710 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 a_10108_32580# VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X711 VDPWR.t44 tdc_0.start_buffer_0.start_delay.t14 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t3 VDPWR.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X712 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t0 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t15 VGND.t553 VGND.t552 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X713 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 VDPWR.t218 VDPWR.t217 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X714 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_1.in.t4 a_25060_11366# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X715 a_24240_21092# variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.out VDPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X716 VGND.t450 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t7 a_16500_15464# VGND.t449 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X717 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t2 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t15 VGND.t492 VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X718 VDPWR.t343 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 VDPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X719 VDPWR.t515 ui_in[4].t6 a_24240_24040# VDPWR.t514 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X720 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 VGND.t167 VGND.t166 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X721 VDPWR.t524 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 VDPWR.t523 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X722 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t319 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X723 VGND.t481 ui_in[1].t0 a_24790_6936# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X724 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 a_10958_32492.t0 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X725 VDPWR.t409 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 VDPWR.t408 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X726 a_16500_11634# VDPWR.t630 VGND.t395 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X727 VDPWR.t587 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 VDPWR.t586 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X728 a_15322_7112# input_stage_0.fine_delay_unit_0.in VDPWR.t475 VDPWR.t474 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X729 VDPWR.t48 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 VDPWR.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X730 a_12420_28316# a_12310_28270# uo_out[2].t2 VDPWR.t136 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X731 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 a_10958_25646.t5 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X732 VGND.t424 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t6 VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X733 a_12420_37822# uo_out[6].t5 VDPWR.t385 VDPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X734 VDPWR.t54 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 VDPWR.t53 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X735 a_25060_14314# ui_in[7].t6 VGND.t296 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X736 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t0 tdc_0.start_buffer_0.start_delay.t15 VGND.t364 VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X737 VGND.t197 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X738 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 VDPWR.t604 VDPWR.t603 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X739 a_10108_32580# tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 a_10958_32492.t5 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X740 variable_delay_dummy_0.out variable_delay_dummy_0.variable_delay_unit_1.in.t5 a_16500_11634# VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X741 a_7140_10670# variable_delay_dummy_0.out VGND.t511 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X742 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 VDPWR.t56 VDPWR.t55 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X743 a_25060_11366# uio_in[0].t6 VGND.t130 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X744 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12308_28732# a_12420_28694# VDPWR.t267 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X745 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 VDPWR.t571 VDPWR.t570 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X746 VDPWR.t582 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 a_12310_39680# VDPWR.t581 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X747 VDPWR.t486 tdc_0.vernier_delay_line_0.stop_strong.t77 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X748 VDPWR.t526 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t13 tdc_0.vernier_delay_line_0.start_neg.t3 VDPWR.t525 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X749 VDPWR.t530 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12420_26034# VDPWR.t529 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X750 a_10958_23364.t11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 a_10108_23452# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X751 a_9330_14924# a_9330_14634# VDPWR.t290 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X752 VDPWR.t358 ui_in[7].t7 a_24240_15196# VDPWR.t357 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X753 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 VGND.t311 VGND.t310 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X754 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 VGND.t530 VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X755 VGND.t451 tdc_0.vernier_delay_line_0.stop_strong.t78 a_10958_39338.t2 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X756 a_13254_39726# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 uo_out[7].t1 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X757 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.start_pos.t14 VDPWR.t595 VDPWR.t594 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X758 input_stage_0.fine_delay_unit_0.in input_stage_0.nand_gate_0.out VGND.t547 VGND.t546 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X759 VDPWR.t424 VDPWR.t422 a_15680_12516# VDPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X760 a_9330_16954.t4 a_9330_15794# VDPWR.t596 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X761 a_10958_32492.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 a_10108_32580# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X762 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 VGND.t520 VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X763 VDPWR.t149 uio_in[0].t7 a_24240_12248# VDPWR.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X764 VGND.t394 VDPWR.t631 a_25060_26106# VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X765 tdc_0.vernier_delay_line_0.stop_strong.t17 a_9330_16954.t36 VDPWR.t28 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X766 tdc_0.vernier_delay_line_0.stop_strong.t16 a_9330_16954.t37 VDPWR.t29 VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X767 tdc_0.vernier_delay_line_0.start_pos.t2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t14 VGND.t14 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X768 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 VGND.t467 VGND.t466 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X769 uo_out[7].t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t102 VDPWR.t101 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X770 VDPWR.t383 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 VDPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X771 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VDPWR.t583 VDPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X772 VGND.t463 ui_in[4].t7 a_25060_23158# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X773 VDPWR.t230 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VDPWR.t229 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X774 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t5 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t14 VDPWR.t591 VDPWR.t590 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X775 VDPWR.t226 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 VDPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X776 a_24240_26988# VDPWR.t419 VDPWR.t421 VDPWR.t420 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X777 a_10108_30826.t4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 a_10958_30210.t5 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X778 VGND.t20 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X779 tdc_0.vernier_delay_line_0.start_neg.t0 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t14 VGND.t128 VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X780 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_5.in.t5 a_24240_23158# VDPWR.t579 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X781 VDPWR.t291 tdc_0.vernier_delay_line_0.stop_strong.t79 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X782 VDPWR.t331 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 VDPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X783 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t511 VDPWR.t510 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X784 VGND.t101 tdc_0.vernier_delay_line_0.start_pos.t15 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X785 a_12420_37444# a_12310_37398# uo_out[6].t2 VDPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X786 VGND.t105 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X787 tdc_0.vernier_delay_line_0.stop_strong.t1 a_9330_16954.t38 VGND.t42 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X788 VGND.t372 tdc_0.start_buffer_0.start_buff.t23 tdc_0.start_buffer_0.start_delay.t0 VGND.t371 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X789 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_4.in.t5 a_24240_20210# VDPWR.t125 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X790 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 VDPWR.t585 VDPWR.t584 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X791 VGND.t437 ui_in[6].t6 a_25060_17262# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X792 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 VDPWR.t247 VDPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X793 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t80 VDPWR.t292 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X794 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 VGND.t319 VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X795 VDPWR.t350 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 VDPWR.t349 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X796 VDPWR.t228 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 a_12310_35116# VDPWR.t227 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X797 VGND.t347 uio_in[2].t0 a_16292_6966# VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X798 VGND.t95 tdc_0.vernier_delay_line_0.stop_strong.t81 a_10958_27928.t6 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X799 VGND.t275 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t2 VGND.t274 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X800 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 VGND.t107 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X801 VDPWR.t389 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12420_35162# VDPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X802 VDPWR.t602 tdc_0.vernier_delay_line_0.start_neg.t14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 VDPWR.t601 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X803 VGND.t7 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t15 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t0 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X804 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 VDPWR.t282 VDPWR.t281 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X805 uo_out[1].t3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t513 VDPWR.t512 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X806 a_25060_17262# ui_in[6].t7 VGND.t438 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X807 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 VGND.t289 VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X808 a_15680_15464# VDPWR.t416 VDPWR.t418 VDPWR.t417 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X809 a_10958_37056.t6 tdc_0.vernier_delay_line_0.stop_strong.t82 VGND.t96 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X810 VDPWR.t362 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 VDPWR.t361 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X811 a_16500_14582# VDPWR.t632 VGND.t392 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X812 VGND.t522 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t15 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t0 VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X813 uo_out[4].t0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 VDPWR.t63 VDPWR.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X814 a_10958_27928.t5 tdc_0.vernier_delay_line_0.stop_strong.t83 VGND.t219 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X815 uo_out[2].t3 a_12310_28270# VGND.t114 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X816 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_1.in.t5 a_24240_11366# VDPWR.t233 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X817 VGND.t383 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 VGND.t382 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X818 VGND.t220 tdc_0.vernier_delay_line_0.stop_strong.t84 a_10958_27928.t4 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X819 a_16500_11634# VDPWR.t633 VGND.t390 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X820 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 VGND.t295 VGND.t294 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X821 a_12420_23752# a_12310_23706# uo_out[0].t1 VDPWR.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X822 VDPWR.t578 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 VDPWR.t577 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X823 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 tdc_0.vernier_delay_line_0.start_neg.t15 VGND.t103 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X824 VGND.t129 tdc_0.vernier_delay_line_0.stop_strong.t85 a_10958_25646.t8 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X825 a_9330_15794# a_9330_15504# VGND.t178 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X826 VGND.t277 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X827 a_13254_28694# uo_out[2].t5 VGND.t283 VGND.t282 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X828 a_10108_39426# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X829 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 tdc_0.vernier_delay_line_0.stop_strong.t86 VDPWR.t145 VDPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X830 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12308_24168# a_12420_24130# VDPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X831 input_stage_1.fine_delay_unit_1.in a_23820_7082# VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X832 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 VGND.t273 VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X833 VDPWR.t532 uio_in[5].t1 input_stage_0.nand_gate_0.out VDPWR.t531 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X834 VDPWR.t283 tdc_0.vernier_delay_line_0.stop_strong.t87 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 VDPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X835 tdc_0.vernier_delay_line_0.stop_strong.t0 a_9330_16954.t39 VGND.t41 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
R0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 552.84
R1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 552.84
R2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 552.84
R3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 552.84
R4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 539.841
R5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 539.841
R6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 539.841
R7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 539.841
R8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 215.293
R9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 215.293
R10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 215.293
R11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 215.293
R12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 166.468
R13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 166.149
R14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 165.8
R15 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 165.8
R16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 85.1574
R17 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 83.8097
R18 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 83.8097
R19 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 83.7172
R20 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 74.288
R21 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 67.7574
R22 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 36.1505
R23 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 36.1505
R24 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 34.5438
R25 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 34.5438
R26 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 17.4005
R27 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 17.4005
R28 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 16.09
R29 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 11.8364
R30 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 9.52217
R31 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 9.52217
R32 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 5.96628
R33 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 5.83219
R34 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 5.74235
R35 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 5.49235
R36 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 1.44072
R37 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 1.32081
R38 VDPWR.n1210 VDPWR.n1209 2207.5
R39 VDPWR.n1226 VDPWR.n1225 2207.5
R40 VDPWR.n1242 VDPWR.n1241 2207.5
R41 VDPWR.n1258 VDPWR.n1257 2207.5
R42 VDPWR.n1274 VDPWR.n1273 2207.5
R43 VDPWR.n1290 VDPWR.n1289 2207.5
R44 VDPWR.n1306 VDPWR.n1305 2207.5
R45 VDPWR.n1322 VDPWR.n1321 2207.5
R46 VDPWR.n1400 VDPWR.n1374 2207.5
R47 VDPWR.n1420 VDPWR.n1374 2207.5
R48 VDPWR.n1422 VDPWR.n1373 2207.5
R49 VDPWR.n1428 VDPWR.n1373 2207.5
R50 VDPWR.n1426 VDPWR.n1358 2207.5
R51 VDPWR.n1448 VDPWR.n1358 2207.5
R52 VDPWR.n1450 VDPWR.n1357 2207.5
R53 VDPWR.n1456 VDPWR.n1357 2207.5
R54 VDPWR.n1454 VDPWR.n1342 2207.5
R55 VDPWR.n1476 VDPWR.n1342 2207.5
R56 VDPWR.n1478 VDPWR.n1341 2207.5
R57 VDPWR.n1007 VDPWR.n1001 2106.47
R58 VDPWR.n1025 VDPWR.n1019 2106.47
R59 VDPWR.n1043 VDPWR.n1037 2106.47
R60 VDPWR.n1061 VDPWR.n1055 2106.47
R61 VDPWR.n1079 VDPWR.n1073 2106.47
R62 VDPWR.n1097 VDPWR.n1091 2106.47
R63 VDPWR.n1115 VDPWR.n1109 2106.47
R64 VDPWR.n1133 VDPWR.n1127 2106.47
R65 VDPWR.n1003 VDPWR.n1002 2101.76
R66 VDPWR.n1021 VDPWR.n1020 2101.76
R67 VDPWR.n1039 VDPWR.n1038 2101.76
R68 VDPWR.n1057 VDPWR.n1056 2101.76
R69 VDPWR.n1075 VDPWR.n1074 2101.76
R70 VDPWR.n1093 VDPWR.n1092 2101.76
R71 VDPWR.n1111 VDPWR.n1110 2101.76
R72 VDPWR.n1129 VDPWR.n1128 2101.76
R73 VDPWR.n1194 VDPWR.n1189 2093.75
R74 VDPWR.n1395 VDPWR.n1389 2093.75
R75 VDPWR.n1199 VDPWR.n1190 2088.75
R76 VDPWR.n1404 VDPWR.n1390 2088.75
R77 VDPWR.n1211 VDPWR.n1209 2070
R78 VDPWR.n1227 VDPWR.n1225 2070
R79 VDPWR.n1243 VDPWR.n1241 2070
R80 VDPWR.n1259 VDPWR.n1257 2070
R81 VDPWR.n1275 VDPWR.n1273 2070
R82 VDPWR.n1291 VDPWR.n1289 2070
R83 VDPWR.n1307 VDPWR.n1305 2070
R84 VDPWR.n1323 VDPWR.n1321 2070
R85 VDPWR.n1480 VDPWR.n1341 2070
R86 VDPWR.n203 VDPWR.n200 1689.71
R87 VDPWR.n469 VDPWR.n200 1689.71
R88 VDPWR.n473 VDPWR.n199 1689.71
R89 VDPWR.n473 VDPWR.n198 1689.71
R90 VDPWR.n227 VDPWR.n224 1689.71
R91 VDPWR.n443 VDPWR.n224 1689.71
R92 VDPWR.n447 VDPWR.n223 1689.71
R93 VDPWR.n447 VDPWR.n222 1689.71
R94 VDPWR.n251 VDPWR.n248 1689.71
R95 VDPWR.n417 VDPWR.n248 1689.71
R96 VDPWR.n421 VDPWR.n247 1689.71
R97 VDPWR.n421 VDPWR.n246 1689.71
R98 VDPWR.n275 VDPWR.n272 1689.71
R99 VDPWR.n391 VDPWR.n272 1689.71
R100 VDPWR.n395 VDPWR.n271 1689.71
R101 VDPWR.n395 VDPWR.n270 1689.71
R102 VDPWR.n299 VDPWR.n296 1689.71
R103 VDPWR.n365 VDPWR.n296 1689.71
R104 VDPWR.n369 VDPWR.n295 1689.71
R105 VDPWR.n369 VDPWR.n294 1689.71
R106 VDPWR.n323 VDPWR.n320 1689.71
R107 VDPWR.n331 VDPWR.n320 1689.71
R108 VDPWR.n335 VDPWR.n319 1689.71
R109 VDPWR.n335 VDPWR.n318 1689.71
R110 VDPWR.n32 VDPWR.n29 1689.71
R111 VDPWR.n98 VDPWR.n29 1689.71
R112 VDPWR.n102 VDPWR.n28 1689.71
R113 VDPWR.n102 VDPWR.n27 1689.71
R114 VDPWR.n56 VDPWR.n53 1689.71
R115 VDPWR.n64 VDPWR.n53 1689.71
R116 VDPWR.n68 VDPWR.n52 1689.71
R117 VDPWR.n68 VDPWR.n51 1689.71
R118 VDPWR.n707 VDPWR.n540 1508.99
R119 VDPWR.n690 VDPWR.n545 1508.99
R120 VDPWR.n673 VDPWR.n550 1508.99
R121 VDPWR.n656 VDPWR.n555 1508.99
R122 VDPWR.n639 VDPWR.n560 1508.99
R123 VDPWR.n622 VDPWR.n565 1508.99
R124 VDPWR.n605 VDPWR.n570 1508.99
R125 VDPWR.n588 VDPWR.n575 1508.99
R126 VDPWR.n1004 VDPWR.n1002 1450
R127 VDPWR.n1022 VDPWR.n1020 1450
R128 VDPWR.n1040 VDPWR.n1038 1450
R129 VDPWR.n1058 VDPWR.n1056 1450
R130 VDPWR.n1076 VDPWR.n1074 1450
R131 VDPWR.n1094 VDPWR.n1092 1450
R132 VDPWR.n1112 VDPWR.n1110 1450
R133 VDPWR.n1130 VDPWR.n1128 1450
R134 VDPWR.n531 VDPWR.n528 1348.04
R135 VDPWR.n1573 VDPWR.n164 1348.04
R136 VDPWR.n1195 VDPWR.n1189 1326.32
R137 VDPWR.n1396 VDPWR.n1389 1326.32
R138 VDPWR.n703 VDPWR.n701 1313.33
R139 VDPWR.n686 VDPWR.n684 1313.33
R140 VDPWR.n669 VDPWR.n667 1313.33
R141 VDPWR.n652 VDPWR.n650 1313.33
R142 VDPWR.n635 VDPWR.n633 1313.33
R143 VDPWR.n618 VDPWR.n616 1313.33
R144 VDPWR.n601 VDPWR.n599 1313.33
R145 VDPWR.n584 VDPWR.n582 1313.33
R146 VDPWR.n1513 VDPWR.n1492 1307.92
R147 VDPWR.n1531 VDPWR.n1524 1307.92
R148 VDPWR.n807 VDPWR.n713 1307.92
R149 VDPWR.n864 VDPWR.n806 1307.92
R150 VDPWR.n517 VDPWR.n516 1307.92
R151 VDPWR.n483 VDPWR.n189 1307.92
R152 VDPWR.n483 VDPWR.n190 1307.92
R153 VDPWR.n485 VDPWR.n187 1307.92
R154 VDPWR.n485 VDPWR.n186 1307.92
R155 VDPWR.n457 VDPWR.n213 1307.92
R156 VDPWR.n457 VDPWR.n214 1307.92
R157 VDPWR.n459 VDPWR.n211 1307.92
R158 VDPWR.n459 VDPWR.n210 1307.92
R159 VDPWR.n431 VDPWR.n237 1307.92
R160 VDPWR.n431 VDPWR.n238 1307.92
R161 VDPWR.n433 VDPWR.n235 1307.92
R162 VDPWR.n433 VDPWR.n234 1307.92
R163 VDPWR.n405 VDPWR.n261 1307.92
R164 VDPWR.n405 VDPWR.n262 1307.92
R165 VDPWR.n407 VDPWR.n259 1307.92
R166 VDPWR.n407 VDPWR.n258 1307.92
R167 VDPWR.n379 VDPWR.n285 1307.92
R168 VDPWR.n379 VDPWR.n286 1307.92
R169 VDPWR.n381 VDPWR.n283 1307.92
R170 VDPWR.n381 VDPWR.n282 1307.92
R171 VDPWR.n345 VDPWR.n309 1307.92
R172 VDPWR.n345 VDPWR.n310 1307.92
R173 VDPWR.n347 VDPWR.n307 1307.92
R174 VDPWR.n347 VDPWR.n306 1307.92
R175 VDPWR.n154 VDPWR.n153 1307.92
R176 VDPWR.n112 VDPWR.n18 1307.92
R177 VDPWR.n112 VDPWR.n19 1307.92
R178 VDPWR.n114 VDPWR.n16 1307.92
R179 VDPWR.n114 VDPWR.n15 1307.92
R180 VDPWR.n80 VDPWR.n39 1307.92
R181 VDPWR.n80 VDPWR.n40 1307.92
R182 VDPWR.n78 VDPWR.n42 1307.92
R183 VDPWR.n78 VDPWR.n43 1307.92
R184 VDPWR.n494 VDPWR.n180 1271.17
R185 VDPWR.n505 VDPWR.n174 1271.17
R186 VDPWR.n131 VDPWR.n9 1271.17
R187 VDPWR.n142 VDPWR.n3 1271.17
R188 VDPWR.n1541 VDPWR.n1512 1126.67
R189 VDPWR.n1515 VDPWR.n1514 1126.67
R190 VDPWR.n1517 VDPWR.n1516 1126.67
R191 VDPWR.n1519 VDPWR.n1518 1126.67
R192 VDPWR.n1521 VDPWR.n1520 1126.67
R193 VDPWR.n1523 VDPWR.n1522 1126.67
R194 VDPWR.n1539 VDPWR.n1526 1126.67
R195 VDPWR.n809 VDPWR.n808 1126.67
R196 VDPWR.n811 VDPWR.n810 1126.67
R197 VDPWR.n813 VDPWR.n812 1126.67
R198 VDPWR.n815 VDPWR.n814 1126.67
R199 VDPWR.n817 VDPWR.n816 1126.67
R200 VDPWR.n819 VDPWR.n818 1126.67
R201 VDPWR.n821 VDPWR.n820 1126.67
R202 VDPWR.n823 VDPWR.n822 1126.67
R203 VDPWR.n825 VDPWR.n824 1126.67
R204 VDPWR.n827 VDPWR.n826 1126.67
R205 VDPWR.n829 VDPWR.n828 1126.67
R206 VDPWR.n831 VDPWR.n830 1126.67
R207 VDPWR.n833 VDPWR.n832 1126.67
R208 VDPWR.n835 VDPWR.n834 1126.67
R209 VDPWR.n837 VDPWR.n836 1126.67
R210 VDPWR.n839 VDPWR.n838 1126.67
R211 VDPWR.n841 VDPWR.n840 1126.67
R212 VDPWR.n843 VDPWR.n842 1126.67
R213 VDPWR.n845 VDPWR.n844 1126.67
R214 VDPWR.n847 VDPWR.n846 1126.67
R215 VDPWR.n849 VDPWR.n848 1126.67
R216 VDPWR.n851 VDPWR.n850 1126.67
R217 VDPWR.n853 VDPWR.n852 1126.67
R218 VDPWR.n855 VDPWR.n854 1126.67
R219 VDPWR.n857 VDPWR.n856 1126.67
R220 VDPWR.n862 VDPWR.n861 1126.67
R221 VDPWR.n859 VDPWR.n858 1126.67
R222 VDPWR.n353 VDPWR.t442 628.097
R223 VDPWR.n120 VDPWR.t437 628.097
R224 VDPWR.n86 VDPWR.t445 628.097
R225 VDPWR.n354 VDPWR.t434 622.766
R226 VDPWR.n121 VDPWR.t422 622.766
R227 VDPWR.n87 VDPWR.t431 622.766
R228 VDPWR.n169 VDPWR.t425 564.04
R229 VDPWR.n519 VDPWR.n516 551.179
R230 VDPWR.n156 VDPWR.n153 551.179
R231 VDPWR.n352 VDPWR.t451 543.053
R232 VDPWR.n119 VDPWR.t428 543.053
R233 VDPWR.n85 VDPWR.t440 543.053
R234 VDPWR.n353 VDPWR.t419 523.774
R235 VDPWR.n120 VDPWR.t448 523.774
R236 VDPWR.n86 VDPWR.t416 523.774
R237 VDPWR.n169 VDPWR.t627 511.623
R238 VDPWR.n531 VDPWR.n530 485.663
R239 VDPWR.n1571 VDPWR.n164 485.663
R240 VDPWR.n484 VDPWR.n188 460.678
R241 VDPWR.n458 VDPWR.n212 460.678
R242 VDPWR.n432 VDPWR.n236 460.678
R243 VDPWR.n406 VDPWR.n260 460.678
R244 VDPWR.n380 VDPWR.n284 460.678
R245 VDPWR.n346 VDPWR.n308 460.678
R246 VDPWR.n113 VDPWR.n17 460.678
R247 VDPWR.n79 VDPWR.n41 460.678
R248 VDPWR.n182 VDPWR.n180 408.981
R249 VDPWR.n176 VDPWR.n174 408.981
R250 VDPWR.n11 VDPWR.n9 408.981
R251 VDPWR.n5 VDPWR.n3 408.981
R252 VDPWR.n706 VDPWR.n699 358.526
R253 VDPWR.n689 VDPWR.n682 358.526
R254 VDPWR.n672 VDPWR.n665 358.526
R255 VDPWR.n655 VDPWR.n648 358.526
R256 VDPWR.n638 VDPWR.n631 358.526
R257 VDPWR.n621 VDPWR.n614 358.526
R258 VDPWR.n604 VDPWR.n597 358.526
R259 VDPWR.n587 VDPWR.n580 358.526
R260 VDPWR.n471 VDPWR.n470 332.803
R261 VDPWR.n445 VDPWR.n444 332.803
R262 VDPWR.n419 VDPWR.n418 332.803
R263 VDPWR.n393 VDPWR.n392 332.803
R264 VDPWR.n367 VDPWR.n366 332.803
R265 VDPWR.n333 VDPWR.n332 332.803
R266 VDPWR.n100 VDPWR.n99 332.803
R267 VDPWR.n66 VDPWR.n65 332.803
R268 VDPWR.n497 VDPWR.n496 313.632
R269 VDPWR.n134 VDPWR.n133 313.632
R270 VDPWR.n508 VDPWR.n507 312.635
R271 VDPWR.n145 VDPWR.n144 312.635
R272 VDPWR.n355 VDPWR.t623 304.647
R273 VDPWR.n355 VDPWR.t629 304.647
R274 VDPWR.n122 VDPWR.t630 304.647
R275 VDPWR.n122 VDPWR.t633 304.647
R276 VDPWR.n88 VDPWR.t625 304.647
R277 VDPWR.n88 VDPWR.t632 304.647
R278 VDPWR.n698 VDPWR.n696 254.195
R279 VDPWR.n681 VDPWR.n679 254.195
R280 VDPWR.n664 VDPWR.n662 254.195
R281 VDPWR.n647 VDPWR.n645 254.195
R282 VDPWR.n630 VDPWR.n628 254.195
R283 VDPWR.n613 VDPWR.n611 254.195
R284 VDPWR.n596 VDPWR.n594 254.195
R285 VDPWR.n579 VDPWR.n577 254.195
R286 VDPWR.n1216 VDPWR.n1208 235.468
R287 VDPWR.n1232 VDPWR.n1224 235.468
R288 VDPWR.n1248 VDPWR.n1240 235.468
R289 VDPWR.n1264 VDPWR.n1256 235.468
R290 VDPWR.n1280 VDPWR.n1272 235.468
R291 VDPWR.n1296 VDPWR.n1288 235.468
R292 VDPWR.n1312 VDPWR.n1304 235.468
R293 VDPWR.n1328 VDPWR.n1320 235.468
R294 VDPWR.n1418 VDPWR.n1379 235.468
R295 VDPWR.n1419 VDPWR.n1418 235.468
R296 VDPWR.n1433 VDPWR.n1372 235.468
R297 VDPWR.n1433 VDPWR.n1367 235.468
R298 VDPWR.n1446 VDPWR.n1363 235.468
R299 VDPWR.n1447 VDPWR.n1446 235.468
R300 VDPWR.n1461 VDPWR.n1356 235.468
R301 VDPWR.n1461 VDPWR.n1351 235.468
R302 VDPWR.n1474 VDPWR.n1347 235.468
R303 VDPWR.n1475 VDPWR.n1474 235.468
R304 VDPWR.n1485 VDPWR.n1340 235.468
R305 VDPWR.n1009 VDPWR.n1000 224.69
R306 VDPWR.n1027 VDPWR.n1018 224.69
R307 VDPWR.n1045 VDPWR.n1036 224.69
R308 VDPWR.n1063 VDPWR.n1054 224.69
R309 VDPWR.n1081 VDPWR.n1072 224.69
R310 VDPWR.n1099 VDPWR.n1090 224.69
R311 VDPWR.n1117 VDPWR.n1108 224.69
R312 VDPWR.n1135 VDPWR.n1126 224.69
R313 VDPWR.n1008 VDPWR.n994 224.189
R314 VDPWR.n1026 VDPWR.n990 224.189
R315 VDPWR.n1044 VDPWR.n986 224.189
R316 VDPWR.n1062 VDPWR.n982 224.189
R317 VDPWR.n1080 VDPWR.n978 224.189
R318 VDPWR.n1098 VDPWR.n974 224.189
R319 VDPWR.n1116 VDPWR.n970 224.189
R320 VDPWR.n1134 VDPWR.n966 224.189
R321 VDPWR.n1193 VDPWR.n1188 223.333
R322 VDPWR.n1394 VDPWR.n1388 223.333
R323 VDPWR.n1200 VDPWR.n1183 222.8
R324 VDPWR.n1405 VDPWR.n1383 222.8
R325 VDPWR.n352 VDPWR.t621 221.72
R326 VDPWR.n119 VDPWR.t626 221.72
R327 VDPWR.n85 VDPWR.t622 221.72
R328 VDPWR.n1216 VDPWR.n1178 220.8
R329 VDPWR.n1232 VDPWR.n1173 220.8
R330 VDPWR.n1248 VDPWR.n1168 220.8
R331 VDPWR.n1264 VDPWR.n1163 220.8
R332 VDPWR.n1280 VDPWR.n1158 220.8
R333 VDPWR.n1296 VDPWR.n1153 220.8
R334 VDPWR.n1312 VDPWR.n1148 220.8
R335 VDPWR.n1328 VDPWR.n1143 220.8
R336 VDPWR.n1485 VDPWR.n1335 220.8
R337 VDPWR.n125 VDPWR.n119 219.549
R338 VDPWR.n91 VDPWR.n85 219.531
R339 VDPWR.n358 VDPWR.n352 219.526
R340 VDPWR.n355 VDPWR.t631 202.44
R341 VDPWR.n122 VDPWR.t628 202.44
R342 VDPWR.n88 VDPWR.t624 202.44
R343 VDPWR.n705 VDPWR.n704 185.162
R344 VDPWR.n688 VDPWR.n687 185.162
R345 VDPWR.n671 VDPWR.n670 185.162
R346 VDPWR.n654 VDPWR.n653 185.162
R347 VDPWR.n637 VDPWR.n636 185.162
R348 VDPWR.n620 VDPWR.n619 185.162
R349 VDPWR.n603 VDPWR.n602 185.162
R350 VDPWR.n586 VDPWR.n585 185.162
R351 VDPWR.n706 VDPWR.n705 185
R352 VDPWR.n689 VDPWR.n688 185
R353 VDPWR.n672 VDPWR.n671 185
R354 VDPWR.n655 VDPWR.n654 185
R355 VDPWR.n638 VDPWR.n637 185
R356 VDPWR.n621 VDPWR.n620 185
R357 VDPWR.n604 VDPWR.n603 185
R358 VDPWR.n587 VDPWR.n586 185
R359 VDPWR.n1514 VDPWR.n1492 181.25
R360 VDPWR.n1514 VDPWR.n1494 181.25
R361 VDPWR.n1516 VDPWR.n1494 181.25
R362 VDPWR.n1516 VDPWR.n1499 181.25
R363 VDPWR.n1518 VDPWR.n1499 181.25
R364 VDPWR.n1518 VDPWR.n1501 181.25
R365 VDPWR.n1520 VDPWR.n1501 181.25
R366 VDPWR.n1520 VDPWR.n1506 181.25
R367 VDPWR.n1522 VDPWR.n1506 181.25
R368 VDPWR.n1522 VDPWR.n1508 181.25
R369 VDPWR.n1512 VDPWR.n1508 181.25
R370 VDPWR.n1529 VDPWR.n1512 181.25
R371 VDPWR.n1529 VDPWR.n1526 181.25
R372 VDPWR.n1531 VDPWR.n1526 181.25
R373 VDPWR.n808 VDPWR.n713 181.25
R374 VDPWR.n808 VDPWR.n715 181.25
R375 VDPWR.n810 VDPWR.n715 181.25
R376 VDPWR.n810 VDPWR.n720 181.25
R377 VDPWR.n812 VDPWR.n720 181.25
R378 VDPWR.n812 VDPWR.n722 181.25
R379 VDPWR.n814 VDPWR.n722 181.25
R380 VDPWR.n814 VDPWR.n727 181.25
R381 VDPWR.n816 VDPWR.n727 181.25
R382 VDPWR.n816 VDPWR.n729 181.25
R383 VDPWR.n818 VDPWR.n729 181.25
R384 VDPWR.n818 VDPWR.n734 181.25
R385 VDPWR.n820 VDPWR.n734 181.25
R386 VDPWR.n820 VDPWR.n736 181.25
R387 VDPWR.n822 VDPWR.n736 181.25
R388 VDPWR.n822 VDPWR.n741 181.25
R389 VDPWR.n824 VDPWR.n741 181.25
R390 VDPWR.n824 VDPWR.n743 181.25
R391 VDPWR.n826 VDPWR.n743 181.25
R392 VDPWR.n826 VDPWR.n748 181.25
R393 VDPWR.n828 VDPWR.n748 181.25
R394 VDPWR.n828 VDPWR.n750 181.25
R395 VDPWR.n830 VDPWR.n750 181.25
R396 VDPWR.n830 VDPWR.n755 181.25
R397 VDPWR.n832 VDPWR.n755 181.25
R398 VDPWR.n832 VDPWR.n757 181.25
R399 VDPWR.n834 VDPWR.n757 181.25
R400 VDPWR.n834 VDPWR.n762 181.25
R401 VDPWR.n836 VDPWR.n762 181.25
R402 VDPWR.n836 VDPWR.n764 181.25
R403 VDPWR.n838 VDPWR.n764 181.25
R404 VDPWR.n838 VDPWR.n769 181.25
R405 VDPWR.n840 VDPWR.n769 181.25
R406 VDPWR.n840 VDPWR.n771 181.25
R407 VDPWR.n842 VDPWR.n771 181.25
R408 VDPWR.n842 VDPWR.n776 181.25
R409 VDPWR.n844 VDPWR.n776 181.25
R410 VDPWR.n844 VDPWR.n778 181.25
R411 VDPWR.n846 VDPWR.n778 181.25
R412 VDPWR.n846 VDPWR.n783 181.25
R413 VDPWR.n848 VDPWR.n783 181.25
R414 VDPWR.n848 VDPWR.n785 181.25
R415 VDPWR.n850 VDPWR.n785 181.25
R416 VDPWR.n850 VDPWR.n790 181.25
R417 VDPWR.n852 VDPWR.n790 181.25
R418 VDPWR.n852 VDPWR.n792 181.25
R419 VDPWR.n854 VDPWR.n792 181.25
R420 VDPWR.n854 VDPWR.n797 181.25
R421 VDPWR.n856 VDPWR.n797 181.25
R422 VDPWR.n856 VDPWR.n799 181.25
R423 VDPWR.n861 VDPWR.n799 181.25
R424 VDPWR.n861 VDPWR.n804 181.25
R425 VDPWR.n858 VDPWR.n804 181.25
R426 VDPWR.n858 VDPWR.n806 181.25
R427 VDPWR.n467 VDPWR.n204 180.236
R428 VDPWR.n468 VDPWR.n467 180.236
R429 VDPWR.n474 VDPWR.n197 180.236
R430 VDPWR.n474 VDPWR.n193 180.236
R431 VDPWR.n441 VDPWR.n228 180.236
R432 VDPWR.n442 VDPWR.n441 180.236
R433 VDPWR.n448 VDPWR.n221 180.236
R434 VDPWR.n448 VDPWR.n217 180.236
R435 VDPWR.n415 VDPWR.n252 180.236
R436 VDPWR.n416 VDPWR.n415 180.236
R437 VDPWR.n422 VDPWR.n245 180.236
R438 VDPWR.n422 VDPWR.n241 180.236
R439 VDPWR.n389 VDPWR.n276 180.236
R440 VDPWR.n390 VDPWR.n389 180.236
R441 VDPWR.n396 VDPWR.n269 180.236
R442 VDPWR.n396 VDPWR.n265 180.236
R443 VDPWR.n363 VDPWR.n300 180.236
R444 VDPWR.n364 VDPWR.n363 180.236
R445 VDPWR.n370 VDPWR.n293 180.236
R446 VDPWR.n370 VDPWR.n289 180.236
R447 VDPWR.n329 VDPWR.n324 180.236
R448 VDPWR.n330 VDPWR.n329 180.236
R449 VDPWR.n336 VDPWR.n317 180.236
R450 VDPWR.n336 VDPWR.n313 180.236
R451 VDPWR.n96 VDPWR.n33 180.236
R452 VDPWR.n97 VDPWR.n96 180.236
R453 VDPWR.n103 VDPWR.n26 180.236
R454 VDPWR.n103 VDPWR.n22 180.236
R455 VDPWR.n62 VDPWR.n57 180.236
R456 VDPWR.n63 VDPWR.n62 180.236
R457 VDPWR.n69 VDPWR.n50 180.236
R458 VDPWR.n69 VDPWR.n46 180.236
R459 VDPWR.n1215 VDPWR.n1214 171.775
R460 VDPWR.n1231 VDPWR.n1230 171.775
R461 VDPWR.n1247 VDPWR.n1246 171.775
R462 VDPWR.n1263 VDPWR.n1262 171.775
R463 VDPWR.n1279 VDPWR.n1278 171.775
R464 VDPWR.n1295 VDPWR.n1294 171.775
R465 VDPWR.n1311 VDPWR.n1310 171.775
R466 VDPWR.n1327 VDPWR.n1326 171.775
R467 VDPWR.n1399 VDPWR.n1380 171.775
R468 VDPWR.n1432 VDPWR.n1431 171.775
R469 VDPWR.n1425 VDPWR.n1364 171.775
R470 VDPWR.n1460 VDPWR.n1459 171.775
R471 VDPWR.n1453 VDPWR.n1348 171.775
R472 VDPWR.n1484 VDPWR.n1483 171.775
R473 VDPWR.t105 VDPWR.n1001 169.983
R474 VDPWR.t234 VDPWR.n1019 169.983
R475 VDPWR.t191 VDPWR.n1037 169.983
R476 VDPWR.t584 VDPWR.n1055 169.983
R477 VDPWR.t154 VDPWR.n1073 169.983
R478 VDPWR.t401 VDPWR.n1091 169.983
R479 VDPWR.t510 VDPWR.n1109 169.983
R480 VDPWR.t40 VDPWR.n1127 169.983
R481 VDPWR VDPWR.n355 169.071
R482 VDPWR VDPWR.n122 169.071
R483 VDPWR VDPWR.n88 169.071
R484 VDPWR VDPWR.n354 166.244
R485 VDPWR VDPWR.n121 166.244
R486 VDPWR VDPWR.n87 166.244
R487 VDPWR.t581 VDPWR.n1003 164.046
R488 VDPWR.t37 VDPWR.n1021 164.046
R489 VDPWR.t227 VDPWR.n1039 164.046
R490 VDPWR.t564 VDPWR.n1057 164.046
R491 VDPWR.t68 VDPWR.n1075 164.046
R492 VDPWR.t337 VDPWR.n1093 164.046
R493 VDPWR.t572 VDPWR.n1111 164.046
R494 VDPWR.t394 VDPWR.n1129 164.046
R495 VDPWR.n203 VDPWR.t477 163.724
R496 VDPWR.t339 VDPWR.n199 163.724
R497 VDPWR.n227 VDPWR.t575 163.724
R498 VDPWR.t502 VDPWR.n223 163.724
R499 VDPWR.n251 VDPWR.t80 163.724
R500 VDPWR.t326 VDPWR.n247 163.724
R501 VDPWR.n275 VDPWR.t552 163.724
R502 VDPWR.t353 VDPWR.n271 163.724
R503 VDPWR.n299 VDPWR.t120 163.724
R504 VDPWR.t204 VDPWR.n295 163.724
R505 VDPWR.n323 VDPWR.t443 163.724
R506 VDPWR.t242 VDPWR.n319 163.724
R507 VDPWR.n32 VDPWR.t438 163.724
R508 VDPWR.t379 VDPWR.n28 163.724
R509 VDPWR.n56 VDPWR.t446 163.724
R510 VDPWR.t484 VDPWR.n52 163.724
R511 VDPWR.n170 VDPWR.n169 161.3
R512 VDPWR.n590 VDPWR.n589 160.959
R513 VDPWR.n607 VDPWR.n606 160.959
R514 VDPWR.n624 VDPWR.n623 160.959
R515 VDPWR.n641 VDPWR.n640 160.959
R516 VDPWR.n658 VDPWR.n657 160.959
R517 VDPWR.n675 VDPWR.n674 160.959
R518 VDPWR.n692 VDPWR.n691 160.959
R519 VDPWR.n709 VDPWR.n708 160.959
R520 VDPWR.n1195 VDPWR.n1188 158.292
R521 VDPWR.n1396 VDPWR.n1388 158.292
R522 VDPWR.n1008 VDPWR.n996 154.667
R523 VDPWR.n1026 VDPWR.n992 154.667
R524 VDPWR.n1044 VDPWR.n988 154.667
R525 VDPWR.n1062 VDPWR.n984 154.667
R526 VDPWR.n1080 VDPWR.n980 154.667
R527 VDPWR.n1098 VDPWR.n976 154.667
R528 VDPWR.n1116 VDPWR.n972 154.667
R529 VDPWR.n1134 VDPWR.n968 154.667
R530 VDPWR.n704 VDPWR.n703 153.304
R531 VDPWR.n687 VDPWR.n686 153.304
R532 VDPWR.n670 VDPWR.n669 153.304
R533 VDPWR.n653 VDPWR.n652 153.304
R534 VDPWR.n636 VDPWR.n635 153.304
R535 VDPWR.n619 VDPWR.n618 153.304
R536 VDPWR.n602 VDPWR.n601 153.304
R537 VDPWR.n585 VDPWR.n584 153.304
R538 VDPWR.t506 VDPWR.n1194 151.868
R539 VDPWR.t550 VDPWR.n1210 151.868
R540 VDPWR.t287 VDPWR.n1226 151.868
R541 VDPWR.t410 VDPWR.n1242 151.868
R542 VDPWR.t182 VDPWR.n1258 151.868
R543 VDPWR.t459 VDPWR.n1274 151.868
R544 VDPWR.t112 VDPWR.n1290 151.868
R545 VDPWR.t55 VDPWR.n1306 151.868
R546 VDPWR.t298 VDPWR.n1322 151.868
R547 VDPWR.t158 VDPWR.n1395 151.868
R548 VDPWR.n1540 VDPWR.n1525 151.03
R549 VDPWR.n470 VDPWR.t39 145.224
R550 VDPWR.t233 VDPWR.n471 145.224
R551 VDPWR.n444 VDPWR.t61 145.224
R552 VDPWR.t516 VDPWR.n445 145.224
R553 VDPWR.n418 VDPWR.t42 145.224
R554 VDPWR.t289 VDPWR.n419 145.224
R555 VDPWR.n392 VDPWR.t473 145.224
R556 VDPWR.t125 VDPWR.n393 145.224
R557 VDPWR.n366 VDPWR.t14 145.224
R558 VDPWR.t579 VDPWR.n367 145.224
R559 VDPWR.n332 VDPWR.t83 145.224
R560 VDPWR.t100 VDPWR.n333 145.224
R561 VDPWR.n99 VDPWR.t548 145.224
R562 VDPWR.t115 VDPWR.n100 145.224
R563 VDPWR.n65 VDPWR.t84 145.224
R564 VDPWR.t606 VDPWR.n66 145.224
R565 VDPWR.n532 VDPWR.n527 143.792
R566 VDPWR.n532 VDPWR.n167 143.792
R567 VDPWR.n1574 VDPWR.n163 143.792
R568 VDPWR.n1570 VDPWR.n163 143.792
R569 VDPWR.n1005 VDPWR.t57 143.49
R570 VDPWR.n1023 VDPWR.t617 143.49
R571 VDPWR.n1041 VDPWR.t388 143.49
R572 VDPWR.n1059 VDPWR.t566 143.49
R573 VDPWR.n1077 VDPWR.t240 143.49
R574 VDPWR.n1095 VDPWR.t134 143.49
R575 VDPWR.n1113 VDPWR.t529 143.49
R576 VDPWR.n1131 VDPWR.t613 143.49
R577 VDPWR.n1006 VDPWR.t272 141.511
R578 VDPWR.n1024 VDPWR.t384 141.511
R579 VDPWR.n1042 VDPWR.t482 141.511
R580 VDPWR.n1060 VDPWR.t588 141.511
R581 VDPWR.n1078 VDPWR.t210 141.511
R582 VDPWR.n1096 VDPWR.t324 141.511
R583 VDPWR.n1114 VDPWR.t294 141.511
R584 VDPWR.n1132 VDPWR.t130 141.511
R585 VDPWR.n1562 VDPWR.n1490 139.512
R586 VDPWR.n1536 VDPWR.n1532 139.512
R587 VDPWR.n963 VDPWR.n711 139.512
R588 VDPWR.n870 VDPWR.n865 139.512
R589 VDPWR.n521 VDPWR.n514 139.512
R590 VDPWR.n521 VDPWR.n520 139.512
R591 VDPWR.n482 VDPWR.n191 139.512
R592 VDPWR.n482 VDPWR.n192 139.512
R593 VDPWR.n486 VDPWR.n185 139.512
R594 VDPWR.n486 VDPWR.n183 139.512
R595 VDPWR.n456 VDPWR.n215 139.512
R596 VDPWR.n456 VDPWR.n216 139.512
R597 VDPWR.n460 VDPWR.n209 139.512
R598 VDPWR.n460 VDPWR.n207 139.512
R599 VDPWR.n430 VDPWR.n239 139.512
R600 VDPWR.n430 VDPWR.n240 139.512
R601 VDPWR.n434 VDPWR.n233 139.512
R602 VDPWR.n434 VDPWR.n231 139.512
R603 VDPWR.n404 VDPWR.n263 139.512
R604 VDPWR.n404 VDPWR.n264 139.512
R605 VDPWR.n408 VDPWR.n257 139.512
R606 VDPWR.n408 VDPWR.n255 139.512
R607 VDPWR.n378 VDPWR.n287 139.512
R608 VDPWR.n378 VDPWR.n288 139.512
R609 VDPWR.n382 VDPWR.n281 139.512
R610 VDPWR.n382 VDPWR.n279 139.512
R611 VDPWR.n344 VDPWR.n311 139.512
R612 VDPWR.n344 VDPWR.n312 139.512
R613 VDPWR.n348 VDPWR.n305 139.512
R614 VDPWR.n348 VDPWR.n303 139.512
R615 VDPWR.n158 VDPWR.n151 139.512
R616 VDPWR.n158 VDPWR.n157 139.512
R617 VDPWR.n111 VDPWR.n20 139.512
R618 VDPWR.n111 VDPWR.n21 139.512
R619 VDPWR.n115 VDPWR.n14 139.512
R620 VDPWR.n115 VDPWR.n12 139.512
R621 VDPWR.n81 VDPWR.n38 139.512
R622 VDPWR.n81 VDPWR.n36 139.512
R623 VDPWR.n77 VDPWR.n45 139.512
R624 VDPWR.n77 VDPWR.n44 139.512
R625 VDPWR.n1196 VDPWR.t349 135.981
R626 VDPWR.n1214 VDPWR.t189 135.981
R627 VDPWR.n1230 VDPWR.t206 135.981
R628 VDPWR.n1246 VDPWR.t577 135.981
R629 VDPWR.n1262 VDPWR.t279 135.981
R630 VDPWR.n1278 VDPWR.t457 135.981
R631 VDPWR.n1294 VDPWR.t369 135.981
R632 VDPWR.n1310 VDPWR.t53 135.981
R633 VDPWR.n1326 VDPWR.t49 135.981
R634 VDPWR.n1397 VDPWR.t517 135.981
R635 VDPWR.t313 VDPWR.n1399 135.981
R636 VDPWR.n1431 VDPWR.t560 135.981
R637 VDPWR.t208 VDPWR.n1425 135.981
R638 VDPWR.n1459 VDPWR.t542 135.981
R639 VDPWR.t72 VDPWR.n1453 135.981
R640 VDPWR.n1483 VDPWR.t250 135.981
R641 VDPWR.n493 VDPWR.n179 135.591
R642 VDPWR.n504 VDPWR.n173 135.591
R643 VDPWR.n130 VDPWR.n8 135.591
R644 VDPWR.n141 VDPWR.n2 135.591
R645 VDPWR.t330 VDPWR.n1197 135.049
R646 VDPWR.t586 VDPWR.n1212 135.049
R647 VDPWR.t30 VDPWR.n1228 135.049
R648 VDPWR.t162 VDPWR.n1244 135.049
R649 VDPWR.t167 VDPWR.n1260 135.049
R650 VDPWR.t359 VDPWR.n1276 135.049
R651 VDPWR.t6 VDPWR.n1292 135.049
R652 VDPWR.t382 VDPWR.n1308 135.049
R653 VDPWR.t132 VDPWR.n1324 135.049
R654 VDPWR.t33 VDPWR.n1402 135.049
R655 VDPWR.n1401 VDPWR.t315 135.049
R656 VDPWR.n1421 VDPWR.t311 135.049
R657 VDPWR.t558 VDPWR.n1423 135.049
R658 VDPWR.t143 VDPWR.n1429 135.049
R659 VDPWR.n1427 VDPWR.t487 135.049
R660 VDPWR.n1449 VDPWR.t471 135.049
R661 VDPWR.t320 VDPWR.n1451 135.049
R662 VDPWR.t519 VDPWR.n1457 135.049
R663 VDPWR.n1455 VDPWR.t128 135.049
R664 VDPWR.n1477 VDPWR.t180 135.049
R665 VDPWR.t252 VDPWR.n1479 135.049
R666 VDPWR.t403 VDPWR.n1481 135.049
R667 VDPWR.n707 VDPWR.n696 134.43
R668 VDPWR.n690 VDPWR.n679 134.43
R669 VDPWR.n673 VDPWR.n662 134.43
R670 VDPWR.n656 VDPWR.n645 134.43
R671 VDPWR.n639 VDPWR.n628 134.43
R672 VDPWR.n622 VDPWR.n611 134.43
R673 VDPWR.n605 VDPWR.n594 134.43
R674 VDPWR.n588 VDPWR.n577 134.43
R675 VDPWR.n1198 VDPWR.t570 132.256
R676 VDPWR.n1213 VDPWR.t66 132.256
R677 VDPWR.n1229 VDPWR.t398 132.256
R678 VDPWR.n1245 VDPWR.t603 132.256
R679 VDPWR.n1261 VDPWR.t86 132.256
R680 VDPWR.n1277 VDPWR.t328 132.256
R681 VDPWR.n1293 VDPWR.t4 132.256
R682 VDPWR.n1309 VDPWR.t231 132.256
R683 VDPWR.n1325 VDPWR.t160 132.256
R684 VDPWR.n1403 VDPWR.t146 132.256
R685 VDPWR.n1398 VDPWR.t307 132.256
R686 VDPWR.n1430 VDPWR.t544 132.256
R687 VDPWR.n1424 VDPWR.t363 132.256
R688 VDPWR.n1458 VDPWR.t494 132.256
R689 VDPWR.n1452 VDPWR.t178 132.256
R690 VDPWR.n1482 VDPWR.t35 132.256
R691 VDPWR.n701 VDPWR.n700 129.874
R692 VDPWR.n700 VDPWR.n696 129.874
R693 VDPWR.n684 VDPWR.n683 129.874
R694 VDPWR.n683 VDPWR.n679 129.874
R695 VDPWR.n667 VDPWR.n666 129.874
R696 VDPWR.n666 VDPWR.n662 129.874
R697 VDPWR.n650 VDPWR.n649 129.874
R698 VDPWR.n649 VDPWR.n645 129.874
R699 VDPWR.n633 VDPWR.n632 129.874
R700 VDPWR.n632 VDPWR.n628 129.874
R701 VDPWR.n616 VDPWR.n615 129.874
R702 VDPWR.n615 VDPWR.n611 129.874
R703 VDPWR.n599 VDPWR.n598 129.874
R704 VDPWR.n598 VDPWR.n594 129.874
R705 VDPWR.n582 VDPWR.n581 129.874
R706 VDPWR.n581 VDPWR.n577 129.874
R707 VDPWR.n498 VDPWR.n177 129.013
R708 VDPWR.n509 VDPWR.n171 129.013
R709 VDPWR.n135 VDPWR.n6 129.013
R710 VDPWR.n146 VDPWR.n0 129.013
R711 VDPWR.n1561 VDPWR.n1493 120.178
R712 VDPWR.n1497 VDPWR.n1495 120.178
R713 VDPWR.n1554 VDPWR.n1500 120.178
R714 VDPWR.n1504 VDPWR.n1502 120.178
R715 VDPWR.n1547 VDPWR.n1507 120.178
R716 VDPWR.n1538 VDPWR.n1537 120.178
R717 VDPWR.n1542 VDPWR.n1509 120.178
R718 VDPWR.n962 VDPWR.n714 120.178
R719 VDPWR.n718 VDPWR.n716 120.178
R720 VDPWR.n955 VDPWR.n721 120.178
R721 VDPWR.n725 VDPWR.n723 120.178
R722 VDPWR.n948 VDPWR.n728 120.178
R723 VDPWR.n732 VDPWR.n730 120.178
R724 VDPWR.n941 VDPWR.n735 120.178
R725 VDPWR.n739 VDPWR.n737 120.178
R726 VDPWR.n934 VDPWR.n742 120.178
R727 VDPWR.n746 VDPWR.n744 120.178
R728 VDPWR.n927 VDPWR.n749 120.178
R729 VDPWR.n753 VDPWR.n751 120.178
R730 VDPWR.n920 VDPWR.n756 120.178
R731 VDPWR.n760 VDPWR.n758 120.178
R732 VDPWR.n913 VDPWR.n763 120.178
R733 VDPWR.n767 VDPWR.n765 120.178
R734 VDPWR.n906 VDPWR.n770 120.178
R735 VDPWR.n774 VDPWR.n772 120.178
R736 VDPWR.n899 VDPWR.n777 120.178
R737 VDPWR.n781 VDPWR.n779 120.178
R738 VDPWR.n892 VDPWR.n784 120.178
R739 VDPWR.n788 VDPWR.n786 120.178
R740 VDPWR.n885 VDPWR.n791 120.178
R741 VDPWR.n795 VDPWR.n793 120.178
R742 VDPWR.n878 VDPWR.n798 120.178
R743 VDPWR.n802 VDPWR.n800 120.178
R744 VDPWR.n871 VDPWR.n805 120.178
R745 VDPWR VDPWR.n1401 108.04
R746 VDPWR.n1423 VDPWR 108.04
R747 VDPWR VDPWR.n1427 108.04
R748 VDPWR.n1451 VDPWR 108.04
R749 VDPWR VDPWR.n1455 108.04
R750 VDPWR.n1479 VDPWR 108.04
R751 VDPWR.t477 VDPWR.t221 88.7478
R752 VDPWR.t148 VDPWR.t39 88.7478
R753 VDPWR.t592 VDPWR.t233 88.7478
R754 VDPWR.t341 VDPWR.t339 88.7478
R755 VDPWR.t575 VDPWR.t265 88.7478
R756 VDPWR.t357 VDPWR.t61 88.7478
R757 VDPWR.t94 VDPWR.t516 88.7478
R758 VDPWR.t405 VDPWR.t502 88.7478
R759 VDPWR.t80 VDPWR.t78 88.7478
R760 VDPWR.t51 VDPWR.t42 88.7478
R761 VDPWR.t258 VDPWR.t289 88.7478
R762 VDPWR.t256 VDPWR.t326 88.7478
R763 VDPWR.t552 VDPWR.t554 88.7478
R764 VDPWR.t274 VDPWR.t473 88.7478
R765 VDPWR.t244 VDPWR.t125 88.7478
R766 VDPWR.t355 VDPWR.t353 88.7478
R767 VDPWR.t120 VDPWR.t123 88.7478
R768 VDPWR.t514 VDPWR.t14 88.7478
R769 VDPWR.t202 VDPWR.t579 88.7478
R770 VDPWR.t412 VDPWR.t204 88.7478
R771 VDPWR.t443 VDPWR.t420 88.7478
R772 VDPWR.t435 VDPWR.t83 88.7478
R773 VDPWR.t508 VDPWR.t100 88.7478
R774 VDPWR.t351 VDPWR.t242 88.7478
R775 VDPWR.t438 VDPWR.t449 88.7478
R776 VDPWR.t423 VDPWR.t548 88.7478
R777 VDPWR.t546 VDPWR.t115 88.7478
R778 VDPWR.t277 VDPWR.t379 88.7478
R779 VDPWR.t446 VDPWR.t417 88.7478
R780 VDPWR.t432 VDPWR.t84 88.7478
R781 VDPWR.t611 VDPWR.t606 88.7478
R782 VDPWR.t609 VDPWR.t484 88.7478
R783 VDPWR.n697 VDPWR.t118 88.2668
R784 VDPWR.n680 VDPWR.t185 88.2668
R785 VDPWR.n663 VDPWR.t169 88.2668
R786 VDPWR.n646 VDPWR.t156 88.2668
R787 VDPWR.n629 VDPWR.t187 88.2668
R788 VDPWR.n612 VDPWR.t214 88.2668
R789 VDPWR.n595 VDPWR.t98 88.2668
R790 VDPWR.n578 VDPWR.t103 88.2668
R791 VDPWR.n699 VDPWR.n697 87.3568
R792 VDPWR.n682 VDPWR.n680 87.3568
R793 VDPWR.n665 VDPWR.n663 87.3568
R794 VDPWR.n648 VDPWR.n646 87.3568
R795 VDPWR.n631 VDPWR.n629 87.3568
R796 VDPWR.n614 VDPWR.n612 87.3568
R797 VDPWR.n597 VDPWR.n595 87.3568
R798 VDPWR.n580 VDPWR.n578 87.3568
R799 VDPWR.t212 VDPWR.t105 87.0838
R800 VDPWR.t600 VDPWR.t212 87.0838
R801 VDPWR.t272 VDPWR.t600 87.0838
R802 VDPWR.t57 VDPWR.t85 87.0838
R803 VDPWR.t85 VDPWR.t101 87.0838
R804 VDPWR.t101 VDPWR.t581 87.0838
R805 VDPWR.t96 VDPWR.t234 87.0838
R806 VDPWR.t397 VDPWR.t96 87.0838
R807 VDPWR.t384 VDPWR.t397 87.0838
R808 VDPWR.t617 VDPWR.t197 87.0838
R809 VDPWR.t197 VDPWR.t619 87.0838
R810 VDPWR.t619 VDPWR.t37 87.0838
R811 VDPWR.t229 VDPWR.t191 87.0838
R812 VDPWR.t82 VDPWR.t229 87.0838
R813 VDPWR.t482 VDPWR.t82 87.0838
R814 VDPWR.t388 VDPWR.t171 87.0838
R815 VDPWR.t171 VDPWR.t346 87.0838
R816 VDPWR.t346 VDPWR.t227 87.0838
R817 VDPWR.t562 VDPWR.t584 87.0838
R818 VDPWR.t476 VDPWR.t562 87.0838
R819 VDPWR.t588 VDPWR.t476 87.0838
R820 VDPWR.t566 VDPWR.t194 87.0838
R821 VDPWR.t194 VDPWR.t62 87.0838
R822 VDPWR.t62 VDPWR.t564 87.0838
R823 VDPWR.t200 VDPWR.t154 87.0838
R824 VDPWR.t173 VDPWR.t200 87.0838
R825 VDPWR.t210 VDPWR.t173 87.0838
R826 VDPWR.t240 VDPWR.t32 87.0838
R827 VDPWR.t32 VDPWR.t538 87.0838
R828 VDPWR.t538 VDPWR.t68 87.0838
R829 VDPWR.t335 VDPWR.t401 87.0838
R830 VDPWR.t267 VDPWR.t335 87.0838
R831 VDPWR.t324 VDPWR.t267 87.0838
R832 VDPWR.t134 VDPWR.t136 87.0838
R833 VDPWR.t136 VDPWR.t536 87.0838
R834 VDPWR.t536 VDPWR.t337 87.0838
R835 VDPWR.t344 VDPWR.t510 87.0838
R836 VDPWR.t264 VDPWR.t344 87.0838
R837 VDPWR.t294 VDPWR.t264 87.0838
R838 VDPWR.t529 VDPWR.t195 87.0838
R839 VDPWR.t195 VDPWR.t512 87.0838
R840 VDPWR.t512 VDPWR.t572 87.0838
R841 VDPWR.t116 VDPWR.t40 87.0838
R842 VDPWR.t196 VDPWR.t116 87.0838
R843 VDPWR.t130 VDPWR.t196 87.0838
R844 VDPWR.t613 VDPWR.t15 87.0838
R845 VDPWR.t15 VDPWR.t317 87.0838
R846 VDPWR.t317 VDPWR.t394 87.0838
R847 VDPWR.n571 VDPWR.t283 85.1439
R848 VDPWR.n566 VDPWR.t396 85.1439
R849 VDPWR.n561 VDPWR.t286 85.1439
R850 VDPWR.n556 VDPWR.t188 85.1439
R851 VDPWR.n551 VDPWR.t486 85.1439
R852 VDPWR.n546 VDPWR.t479 85.1439
R853 VDPWR.n541 VDPWR.t216 85.1439
R854 VDPWR.n536 VDPWR.t291 85.1439
R855 VDPWR.n997 VDPWR.t273 85.0216
R856 VDPWR.n1012 VDPWR.t58 85.0216
R857 VDPWR.n993 VDPWR.t385 85.0216
R858 VDPWR.n1030 VDPWR.t618 85.0216
R859 VDPWR.n989 VDPWR.t483 85.0216
R860 VDPWR.n1048 VDPWR.t389 85.0216
R861 VDPWR.n985 VDPWR.t589 85.0216
R862 VDPWR.n1066 VDPWR.t567 85.0216
R863 VDPWR.n981 VDPWR.t211 85.0216
R864 VDPWR.n1084 VDPWR.t241 85.0216
R865 VDPWR.n977 VDPWR.t325 85.0216
R866 VDPWR.n1102 VDPWR.t135 85.0216
R867 VDPWR.n973 VDPWR.t295 85.0216
R868 VDPWR.n1120 VDPWR.t530 85.0216
R869 VDPWR.n969 VDPWR.t131 85.0216
R870 VDPWR.n1138 VDPWR.t614 85.0216
R871 VDPWR.n166 VDPWR.t535 84.9265
R872 VDPWR.n162 VDPWR.t532 84.9265
R873 VDPWR.n1534 VDPWR.t568 84.9238
R874 VDPWR.n1527 VDPWR.t303 84.9238
R875 VDPWR.n48 VDPWR.n47 84.8474
R876 VDPWR.n1491 VDPWR.t284 84.7934
R877 VDPWR.n1558 VDPWR.t172 84.7934
R878 VDPWR.n1498 VDPWR.t89 84.7934
R879 VDPWR.n1551 VDPWR.t302 84.7934
R880 VDPWR.n1505 VDPWR.t304 84.7934
R881 VDPWR.n1544 VDPWR.t301 84.7934
R882 VDPWR.n712 VDPWR.t107 84.7934
R883 VDPWR.n959 VDPWR.t19 84.7934
R884 VDPWR.n719 VDPWR.t25 84.7934
R885 VDPWR.n952 VDPWR.t27 84.7934
R886 VDPWR.n726 VDPWR.t22 84.7934
R887 VDPWR.n945 VDPWR.t21 84.7934
R888 VDPWR.n733 VDPWR.t109 84.7934
R889 VDPWR.n938 VDPWR.t111 84.7934
R890 VDPWR.n740 VDPWR.t24 84.7934
R891 VDPWR.n931 VDPWR.t29 84.7934
R892 VDPWR.n747 VDPWR.t23 84.7934
R893 VDPWR.n924 VDPWR.t28 84.7934
R894 VDPWR.n754 VDPWR.t20 84.7934
R895 VDPWR.n917 VDPWR.t108 84.7934
R896 VDPWR.n761 VDPWR.t110 84.7934
R897 VDPWR.n910 VDPWR.t26 84.7934
R898 VDPWR.n768 VDPWR.t596 84.7934
R899 VDPWR.n903 VDPWR.t598 84.7934
R900 VDPWR.n775 VDPWR.t599 84.7934
R901 VDPWR.n896 VDPWR.t597 84.7934
R902 VDPWR.n782 VDPWR.t193 84.7934
R903 VDPWR.n889 VDPWR.t400 84.7934
R904 VDPWR.n789 VDPWR.t225 84.7934
R905 VDPWR.n882 VDPWR.t290 84.7934
R906 VDPWR.n796 VDPWR.t164 84.7934
R907 VDPWR.n875 VDPWR.t198 84.7934
R908 VDPWR.n803 VDPWR.t574 84.7934
R909 VDPWR.n868 VDPWR.t605 84.7934
R910 VDPWR.n515 VDPWR.t153 84.7934
R911 VDPWR.n480 VDPWR.t300 84.7934
R912 VDPWR.n488 VDPWR.t151 84.7934
R913 VDPWR.n454 VDPWR.t528 84.7934
R914 VDPWR.n462 VDPWR.t533 84.7934
R915 VDPWR.n428 VDPWR.t549 84.7934
R916 VDPWR.n436 VDPWR.t306 84.7934
R917 VDPWR.n402 VDPWR.t75 84.7934
R918 VDPWR.n410 VDPWR.t184 84.7934
R919 VDPWR.n376 VDPWR.t71 84.7934
R920 VDPWR.n384 VDPWR.t122 84.7934
R921 VDPWR.n342 VDPWR.t255 84.7934
R922 VDPWR.n350 VDPWR.t452 84.7934
R923 VDPWR.n152 VDPWR.t608 84.7934
R924 VDPWR.n109 VDPWR.t569 84.7934
R925 VDPWR.n117 VDPWR.t430 84.7934
R926 VDPWR.n75 VDPWR.t138 84.7934
R927 VDPWR.n83 VDPWR.t441 84.7934
R928 VDPWR.n573 VDPWR.t114 84.7906
R929 VDPWR.n571 VDPWR.t104 84.7906
R930 VDPWR.n572 VDPWR.t580 84.7906
R931 VDPWR.n568 VDPWR.t292 84.7906
R932 VDPWR.n566 VDPWR.t293 84.7906
R933 VDPWR.n567 VDPWR.t99 84.7906
R934 VDPWR.n563 VDPWR.t215 84.7906
R935 VDPWR.n561 VDPWR.t348 84.7906
R936 VDPWR.n562 VDPWR.t226 84.7906
R937 VDPWR.n558 VDPWR.t381 84.7906
R938 VDPWR.n556 VDPWR.t583 84.7906
R939 VDPWR.n557 VDPWR.t276 84.7906
R940 VDPWR.n553 VDPWR.t493 84.7906
R941 VDPWR.n551 VDPWR.t157 84.7906
R942 VDPWR.n552 VDPWR.t199 84.7906
R943 VDPWR.n548 VDPWR.t285 84.7906
R944 VDPWR.n546 VDPWR.t170 84.7906
R945 VDPWR.n547 VDPWR.t334 84.7906
R946 VDPWR.n543 VDPWR.t186 84.7906
R947 VDPWR.n541 VDPWR.t407 84.7906
R948 VDPWR.n542 VDPWR.t343 84.7906
R949 VDPWR.n538 VDPWR.t145 84.7906
R950 VDPWR.n536 VDPWR.t319 84.7906
R951 VDPWR.n537 VDPWR.t119 84.7906
R952 VDPWR.n168 VDPWR.t427 84.7879
R953 VDPWR.n534 VDPWR.t534 84.7879
R954 VDPWR.n491 VDPWR.t77 84.7771
R955 VDPWR.n502 VDPWR.t3 84.7771
R956 VDPWR.n128 VDPWR.t166 84.7771
R957 VDPWR.n139 VDPWR.t415 84.7771
R958 VDPWR.n206 VDPWR.n205 84.7744
R959 VDPWR.n195 VDPWR.n194 84.7744
R960 VDPWR.n230 VDPWR.n229 84.7744
R961 VDPWR.n219 VDPWR.n218 84.7744
R962 VDPWR.n254 VDPWR.n253 84.7744
R963 VDPWR.n243 VDPWR.n242 84.7744
R964 VDPWR.n278 VDPWR.n277 84.7744
R965 VDPWR.n267 VDPWR.n266 84.7744
R966 VDPWR.n302 VDPWR.n301 84.7744
R967 VDPWR.n291 VDPWR.n290 84.7744
R968 VDPWR.n326 VDPWR.n325 84.7744
R969 VDPWR.n315 VDPWR.n314 84.7744
R970 VDPWR.n35 VDPWR.n34 84.7744
R971 VDPWR.n24 VDPWR.n23 84.7744
R972 VDPWR.n59 VDPWR.n58 84.7744
R973 VDPWR.n500 VDPWR.t17 84.7716
R974 VDPWR.n511 VDPWR.t462 84.7716
R975 VDPWR.n137 VDPWR.t1 84.7716
R976 VDPWR.n148 VDPWR.t475 84.7716
R977 VDPWR.n206 VDPWR.t478 83.8097
R978 VDPWR.n195 VDPWR.t340 83.8097
R979 VDPWR.n230 VDPWR.t576 83.8097
R980 VDPWR.n219 VDPWR.t503 83.8097
R981 VDPWR.n254 VDPWR.t81 83.8097
R982 VDPWR.n243 VDPWR.t327 83.8097
R983 VDPWR.n278 VDPWR.t553 83.8097
R984 VDPWR.n267 VDPWR.t354 83.8097
R985 VDPWR.n302 VDPWR.t121 83.8097
R986 VDPWR.n291 VDPWR.t205 83.8097
R987 VDPWR.n326 VDPWR.t444 83.8097
R988 VDPWR.n315 VDPWR.t243 83.8097
R989 VDPWR.n35 VDPWR.t439 83.8097
R990 VDPWR.n24 VDPWR.t380 83.8097
R991 VDPWR.n59 VDPWR.t447 83.8097
R992 VDPWR.n48 VDPWR.t485 83.8097
R993 VDPWR.t465 VDPWR.t506 81.9613
R994 VDPWR.t392 VDPWR.t465 81.9613
R995 VDPWR.t349 VDPWR.t392 81.9613
R996 VDPWR.t570 VDPWR.t268 81.9613
R997 VDPWR.t268 VDPWR.t332 81.9613
R998 VDPWR.t332 VDPWR.t330 81.9613
R999 VDPWR.t176 VDPWR.t550 81.9613
R1000 VDPWR.t174 VDPWR.t176 81.9613
R1001 VDPWR.t189 VDPWR.t174 81.9613
R1002 VDPWR.t66 VDPWR.t64 81.9613
R1003 VDPWR.t64 VDPWR.t540 81.9613
R1004 VDPWR.t540 VDPWR.t586 81.9613
R1005 VDPWR.t296 VDPWR.t287 81.9613
R1006 VDPWR.t217 VDPWR.t296 81.9613
R1007 VDPWR.t206 VDPWR.t217 81.9613
R1008 VDPWR.t398 VDPWR.t523 81.9613
R1009 VDPWR.t523 VDPWR.t521 81.9613
R1010 VDPWR.t521 VDPWR.t30 81.9613
R1011 VDPWR.t47 VDPWR.t410 81.9613
R1012 VDPWR.t92 VDPWR.t47 81.9613
R1013 VDPWR.t577 VDPWR.t92 81.9613
R1014 VDPWR.t603 VDPWR.t59 81.9613
R1015 VDPWR.t59 VDPWR.t390 81.9613
R1016 VDPWR.t390 VDPWR.t162 81.9613
R1017 VDPWR.t480 VDPWR.t182 81.9613
R1018 VDPWR.t281 VDPWR.t480 81.9613
R1019 VDPWR.t279 VDPWR.t281 81.9613
R1020 VDPWR.t86 VDPWR.t498 81.9613
R1021 VDPWR.t498 VDPWR.t246 81.9613
R1022 VDPWR.t246 VDPWR.t167 81.9613
R1023 VDPWR.t453 VDPWR.t459 81.9613
R1024 VDPWR.t455 VDPWR.t453 81.9613
R1025 VDPWR.t457 VDPWR.t455 81.9613
R1026 VDPWR.t328 VDPWR.t361 81.9613
R1027 VDPWR.t361 VDPWR.t377 81.9613
R1028 VDPWR.t377 VDPWR.t359 81.9613
R1029 VDPWR.t408 VDPWR.t112 81.9613
R1030 VDPWR.t371 VDPWR.t408 81.9613
R1031 VDPWR.t369 VDPWR.t371 81.9613
R1032 VDPWR.t4 VDPWR.t238 81.9613
R1033 VDPWR.t238 VDPWR.t12 81.9613
R1034 VDPWR.t12 VDPWR.t6 81.9613
R1035 VDPWR.t504 VDPWR.t55 81.9613
R1036 VDPWR.t126 VDPWR.t504 81.9613
R1037 VDPWR.t53 VDPWR.t126 81.9613
R1038 VDPWR.t231 VDPWR.t491 81.9613
R1039 VDPWR.t491 VDPWR.t489 81.9613
R1040 VDPWR.t489 VDPWR.t382 81.9613
R1041 VDPWR.t262 VDPWR.t298 81.9613
R1042 VDPWR.t594 VDPWR.t262 81.9613
R1043 VDPWR.t49 VDPWR.t594 81.9613
R1044 VDPWR.t160 VDPWR.t601 81.9613
R1045 VDPWR.t601 VDPWR.t223 81.9613
R1046 VDPWR.t223 VDPWR.t132 81.9613
R1047 VDPWR.t525 VDPWR.t158 81.9613
R1048 VDPWR.t375 VDPWR.t525 81.9613
R1049 VDPWR.t517 VDPWR.t375 81.9613
R1050 VDPWR.t146 VDPWR.t10 81.9613
R1051 VDPWR.t10 VDPWR.t8 81.9613
R1052 VDPWR.t8 VDPWR.t33 81.9613
R1053 VDPWR.t315 VDPWR.t141 81.9613
R1054 VDPWR.t141 VDPWR.t590 81.9613
R1055 VDPWR.t590 VDPWR.t313 81.9613
R1056 VDPWR.t307 VDPWR.t309 81.9613
R1057 VDPWR.t309 VDPWR.t496 81.9613
R1058 VDPWR.t496 VDPWR.t311 81.9613
R1059 VDPWR.t556 VDPWR.t558 81.9613
R1060 VDPWR.t260 VDPWR.t556 81.9613
R1061 VDPWR.t560 VDPWR.t260 81.9613
R1062 VDPWR.t544 VDPWR.t322 81.9613
R1063 VDPWR.t322 VDPWR.t386 81.9613
R1064 VDPWR.t386 VDPWR.t143 81.9613
R1065 VDPWR.t487 VDPWR.t463 81.9613
R1066 VDPWR.t463 VDPWR.t236 81.9613
R1067 VDPWR.t236 VDPWR.t208 81.9613
R1068 VDPWR.t363 VDPWR.t367 81.9613
R1069 VDPWR.t367 VDPWR.t365 81.9613
R1070 VDPWR.t365 VDPWR.t471 81.9613
R1071 VDPWR.t139 VDPWR.t320 81.9613
R1072 VDPWR.t373 VDPWR.t139 81.9613
R1073 VDPWR.t542 VDPWR.t373 81.9613
R1074 VDPWR.t494 VDPWR.t615 81.9613
R1075 VDPWR.t615 VDPWR.t219 81.9613
R1076 VDPWR.t219 VDPWR.t519 81.9613
R1077 VDPWR.t128 VDPWR.t270 81.9613
R1078 VDPWR.t270 VDPWR.t500 81.9613
R1079 VDPWR.t500 VDPWR.t72 81.9613
R1080 VDPWR.t178 VDPWR.t469 81.9613
R1081 VDPWR.t469 VDPWR.t467 81.9613
R1082 VDPWR.t467 VDPWR.t180 81.9613
R1083 VDPWR.t90 VDPWR.t252 81.9613
R1084 VDPWR.t248 VDPWR.t90 81.9613
R1085 VDPWR.t250 VDPWR.t248 81.9613
R1086 VDPWR.t35 VDPWR.t43 81.9613
R1087 VDPWR.t43 VDPWR.t45 81.9613
R1088 VDPWR.t45 VDPWR.t403 81.9613
R1089 VDPWR.n1392 VDPWR.n1391 75.8478
R1090 VDPWR.n1387 VDPWR.n1386 75.7173
R1091 VDPWR.n1407 VDPWR.n1385 75.7173
R1092 VDPWR.n1408 VDPWR.n1384 75.7173
R1093 VDPWR.n1411 VDPWR.n1382 75.7173
R1094 VDPWR.n1412 VDPWR.n1381 75.7173
R1095 VDPWR.n1416 VDPWR.n1413 75.7173
R1096 VDPWR.n1415 VDPWR.n1414 75.7173
R1097 VDPWR.n1376 VDPWR.n1375 75.7173
R1098 VDPWR.n1371 VDPWR.n1370 75.7173
R1099 VDPWR.n1435 VDPWR.n1369 75.7173
R1100 VDPWR.n1436 VDPWR.n1368 75.7173
R1101 VDPWR.n1439 VDPWR.n1366 75.7173
R1102 VDPWR.n1440 VDPWR.n1365 75.7173
R1103 VDPWR.n1444 VDPWR.n1441 75.7173
R1104 VDPWR.n1443 VDPWR.n1442 75.7173
R1105 VDPWR.n1360 VDPWR.n1359 75.7173
R1106 VDPWR.n1355 VDPWR.n1354 75.7173
R1107 VDPWR.n1463 VDPWR.n1353 75.7173
R1108 VDPWR.n1464 VDPWR.n1352 75.7173
R1109 VDPWR.n1467 VDPWR.n1350 75.7173
R1110 VDPWR.n1468 VDPWR.n1349 75.7173
R1111 VDPWR.n1472 VDPWR.n1469 75.7173
R1112 VDPWR.n1471 VDPWR.n1470 75.7173
R1113 VDPWR.n1344 VDPWR.n1343 75.7173
R1114 VDPWR.n1339 VDPWR.n1338 75.7173
R1115 VDPWR.n1487 VDPWR.n1337 75.7173
R1116 VDPWR.n1488 VDPWR.n1336 75.7173
R1117 VDPWR.n1192 VDPWR.n1191 75.7173
R1118 VDPWR.n1187 VDPWR.n1186 75.7173
R1119 VDPWR.n1202 VDPWR.n1185 75.7173
R1120 VDPWR.n1203 VDPWR.n1184 75.7173
R1121 VDPWR.n1206 VDPWR.n1205 75.7173
R1122 VDPWR.n1182 VDPWR.n1181 75.7173
R1123 VDPWR.n1218 VDPWR.n1180 75.7173
R1124 VDPWR.n1219 VDPWR.n1179 75.7173
R1125 VDPWR.n1222 VDPWR.n1221 75.7173
R1126 VDPWR.n1177 VDPWR.n1176 75.7173
R1127 VDPWR.n1234 VDPWR.n1175 75.7173
R1128 VDPWR.n1235 VDPWR.n1174 75.7173
R1129 VDPWR.n1238 VDPWR.n1237 75.7173
R1130 VDPWR.n1172 VDPWR.n1171 75.7173
R1131 VDPWR.n1250 VDPWR.n1170 75.7173
R1132 VDPWR.n1251 VDPWR.n1169 75.7173
R1133 VDPWR.n1254 VDPWR.n1253 75.7173
R1134 VDPWR.n1167 VDPWR.n1166 75.7173
R1135 VDPWR.n1266 VDPWR.n1165 75.7173
R1136 VDPWR.n1267 VDPWR.n1164 75.7173
R1137 VDPWR.n1270 VDPWR.n1269 75.7173
R1138 VDPWR.n1162 VDPWR.n1161 75.7173
R1139 VDPWR.n1282 VDPWR.n1160 75.7173
R1140 VDPWR.n1283 VDPWR.n1159 75.7173
R1141 VDPWR.n1286 VDPWR.n1285 75.7173
R1142 VDPWR.n1157 VDPWR.n1156 75.7173
R1143 VDPWR.n1298 VDPWR.n1155 75.7173
R1144 VDPWR.n1299 VDPWR.n1154 75.7173
R1145 VDPWR.n1302 VDPWR.n1301 75.7173
R1146 VDPWR.n1152 VDPWR.n1151 75.7173
R1147 VDPWR.n1314 VDPWR.n1150 75.7173
R1148 VDPWR.n1315 VDPWR.n1149 75.7173
R1149 VDPWR.n1318 VDPWR.n1317 75.7173
R1150 VDPWR.n1147 VDPWR.n1146 75.7173
R1151 VDPWR.n1330 VDPWR.n1145 75.7173
R1152 VDPWR.n1331 VDPWR.n1144 75.7173
R1153 VDPWR.n999 VDPWR.n998 75.5
R1154 VDPWR.n1013 VDPWR.n995 75.5
R1155 VDPWR.n1016 VDPWR.n1015 75.5
R1156 VDPWR.n1031 VDPWR.n991 75.5
R1157 VDPWR.n1034 VDPWR.n1033 75.5
R1158 VDPWR.n1049 VDPWR.n987 75.5
R1159 VDPWR.n1052 VDPWR.n1051 75.5
R1160 VDPWR.n1067 VDPWR.n983 75.5
R1161 VDPWR.n1070 VDPWR.n1069 75.5
R1162 VDPWR.n1085 VDPWR.n979 75.5
R1163 VDPWR.n1088 VDPWR.n1087 75.5
R1164 VDPWR.n1103 VDPWR.n975 75.5
R1165 VDPWR.n1106 VDPWR.n1105 75.5
R1166 VDPWR.n1121 VDPWR.n971 75.5
R1167 VDPWR.n1124 VDPWR.n1123 75.5
R1168 VDPWR.n1139 VDPWR.n967 75.5
R1169 VDPWR.n497 VDPWR.n180 61.6672
R1170 VDPWR.n508 VDPWR.n174 61.6672
R1171 VDPWR.n134 VDPWR.n9 61.6672
R1172 VDPWR.n145 VDPWR.n3 61.6672
R1173 VDPWR.n518 VDPWR.t152 57.2869
R1174 VDPWR.n155 VDPWR.t607 57.2869
R1175 VDPWR.n1197 VDPWR 50.2946
R1176 VDPWR.n1212 VDPWR 50.2946
R1177 VDPWR.n1228 VDPWR 50.2946
R1178 VDPWR.n1244 VDPWR 50.2946
R1179 VDPWR.n1260 VDPWR 50.2946
R1180 VDPWR.n1276 VDPWR 50.2946
R1181 VDPWR.n1292 VDPWR 50.2946
R1182 VDPWR.n1308 VDPWR 50.2946
R1183 VDPWR.n1324 VDPWR 50.2946
R1184 VDPWR.n1402 VDPWR 50.2946
R1185 VDPWR VDPWR.n1421 50.2946
R1186 VDPWR.n1429 VDPWR 50.2946
R1187 VDPWR VDPWR.n1449 50.2946
R1188 VDPWR.n1457 VDPWR 50.2946
R1189 VDPWR VDPWR.n1477 50.2946
R1190 VDPWR.n1481 VDPWR 50.2946
R1191 VDPWR.n1536 VDPWR.n1531 46.2505
R1192 VDPWR.n1531 VDPWR.n1525 46.2505
R1193 VDPWR.n1530 VDPWR.n1529 46.2505
R1194 VDPWR.n1529 VDPWR.n1525 46.2505
R1195 VDPWR.n1546 VDPWR.n1508 46.2505
R1196 VDPWR.n1525 VDPWR.n1508 46.2505
R1197 VDPWR.n1548 VDPWR.n1506 46.2505
R1198 VDPWR.n1525 VDPWR.n1506 46.2505
R1199 VDPWR.n1553 VDPWR.n1501 46.2505
R1200 VDPWR.n1525 VDPWR.n1501 46.2505
R1201 VDPWR.n1555 VDPWR.n1499 46.2505
R1202 VDPWR.n1525 VDPWR.n1499 46.2505
R1203 VDPWR.n1560 VDPWR.n1494 46.2505
R1204 VDPWR.n1525 VDPWR.n1494 46.2505
R1205 VDPWR.n1562 VDPWR.n1492 46.2505
R1206 VDPWR.n1525 VDPWR.n1492 46.2505
R1207 VDPWR.n870 VDPWR.n806 46.2505
R1208 VDPWR.n860 VDPWR.n806 46.2505
R1209 VDPWR.n872 VDPWR.n804 46.2505
R1210 VDPWR.n860 VDPWR.n804 46.2505
R1211 VDPWR.n877 VDPWR.n799 46.2505
R1212 VDPWR.n860 VDPWR.n799 46.2505
R1213 VDPWR.n879 VDPWR.n797 46.2505
R1214 VDPWR.n860 VDPWR.n797 46.2505
R1215 VDPWR.n884 VDPWR.n792 46.2505
R1216 VDPWR.n860 VDPWR.n792 46.2505
R1217 VDPWR.n886 VDPWR.n790 46.2505
R1218 VDPWR.n860 VDPWR.n790 46.2505
R1219 VDPWR.n891 VDPWR.n785 46.2505
R1220 VDPWR.n860 VDPWR.n785 46.2505
R1221 VDPWR.n893 VDPWR.n783 46.2505
R1222 VDPWR.n860 VDPWR.n783 46.2505
R1223 VDPWR.n898 VDPWR.n778 46.2505
R1224 VDPWR.n860 VDPWR.n778 46.2505
R1225 VDPWR.n900 VDPWR.n776 46.2505
R1226 VDPWR.n860 VDPWR.n776 46.2505
R1227 VDPWR.n905 VDPWR.n771 46.2505
R1228 VDPWR.n860 VDPWR.n771 46.2505
R1229 VDPWR.n907 VDPWR.n769 46.2505
R1230 VDPWR.n860 VDPWR.n769 46.2505
R1231 VDPWR.n912 VDPWR.n764 46.2505
R1232 VDPWR.n860 VDPWR.n764 46.2505
R1233 VDPWR.n914 VDPWR.n762 46.2505
R1234 VDPWR.n860 VDPWR.n762 46.2505
R1235 VDPWR.n919 VDPWR.n757 46.2505
R1236 VDPWR.n860 VDPWR.n757 46.2505
R1237 VDPWR.n921 VDPWR.n755 46.2505
R1238 VDPWR.n860 VDPWR.n755 46.2505
R1239 VDPWR.n926 VDPWR.n750 46.2505
R1240 VDPWR.n860 VDPWR.n750 46.2505
R1241 VDPWR.n928 VDPWR.n748 46.2505
R1242 VDPWR.n860 VDPWR.n748 46.2505
R1243 VDPWR.n933 VDPWR.n743 46.2505
R1244 VDPWR.n860 VDPWR.n743 46.2505
R1245 VDPWR.n935 VDPWR.n741 46.2505
R1246 VDPWR.n860 VDPWR.n741 46.2505
R1247 VDPWR.n940 VDPWR.n736 46.2505
R1248 VDPWR.n860 VDPWR.n736 46.2505
R1249 VDPWR.n942 VDPWR.n734 46.2505
R1250 VDPWR.n860 VDPWR.n734 46.2505
R1251 VDPWR.n947 VDPWR.n729 46.2505
R1252 VDPWR.n860 VDPWR.n729 46.2505
R1253 VDPWR.n949 VDPWR.n727 46.2505
R1254 VDPWR.n860 VDPWR.n727 46.2505
R1255 VDPWR.n954 VDPWR.n722 46.2505
R1256 VDPWR.n860 VDPWR.n722 46.2505
R1257 VDPWR.n956 VDPWR.n720 46.2505
R1258 VDPWR.n860 VDPWR.n720 46.2505
R1259 VDPWR.n961 VDPWR.n715 46.2505
R1260 VDPWR.n860 VDPWR.n715 46.2505
R1261 VDPWR.n963 VDPWR.n713 46.2505
R1262 VDPWR.n860 VDPWR.n713 46.2505
R1263 VDPWR.n521 VDPWR.n516 46.2505
R1264 VDPWR.n483 VDPWR.n482 46.2505
R1265 VDPWR.n484 VDPWR.n483 46.2505
R1266 VDPWR.n486 VDPWR.n485 46.2505
R1267 VDPWR.n485 VDPWR.n484 46.2505
R1268 VDPWR.n457 VDPWR.n456 46.2505
R1269 VDPWR.n458 VDPWR.n457 46.2505
R1270 VDPWR.n460 VDPWR.n459 46.2505
R1271 VDPWR.n459 VDPWR.n458 46.2505
R1272 VDPWR.n431 VDPWR.n430 46.2505
R1273 VDPWR.n432 VDPWR.n431 46.2505
R1274 VDPWR.n434 VDPWR.n433 46.2505
R1275 VDPWR.n433 VDPWR.n432 46.2505
R1276 VDPWR.n405 VDPWR.n404 46.2505
R1277 VDPWR.n406 VDPWR.n405 46.2505
R1278 VDPWR.n408 VDPWR.n407 46.2505
R1279 VDPWR.n407 VDPWR.n406 46.2505
R1280 VDPWR.n379 VDPWR.n378 46.2505
R1281 VDPWR.n380 VDPWR.n379 46.2505
R1282 VDPWR.n382 VDPWR.n381 46.2505
R1283 VDPWR.n381 VDPWR.n380 46.2505
R1284 VDPWR.n345 VDPWR.n344 46.2505
R1285 VDPWR.n346 VDPWR.n345 46.2505
R1286 VDPWR.n348 VDPWR.n347 46.2505
R1287 VDPWR.n347 VDPWR.n346 46.2505
R1288 VDPWR.n158 VDPWR.n153 46.2505
R1289 VDPWR.n112 VDPWR.n111 46.2505
R1290 VDPWR.n113 VDPWR.n112 46.2505
R1291 VDPWR.n115 VDPWR.n114 46.2505
R1292 VDPWR.n114 VDPWR.n113 46.2505
R1293 VDPWR.n81 VDPWR.n80 46.2505
R1294 VDPWR.n80 VDPWR.n79 46.2505
R1295 VDPWR.n78 VDPWR.n77 46.2505
R1296 VDPWR.n79 VDPWR.n78 46.2505
R1297 VDPWR.n529 VDPWR.t426 44.5923
R1298 VDPWR.n1572 VDPWR.t531 44.5923
R1299 VDPWR.n863 VDPWR.n860 44.5678
R1300 VDPWR.t221 VDPWR.n202 44.3742
R1301 VDPWR.n202 VDPWR.t148 44.3742
R1302 VDPWR.n472 VDPWR.t592 44.3742
R1303 VDPWR.n472 VDPWR.t341 44.3742
R1304 VDPWR.t265 VDPWR.n226 44.3742
R1305 VDPWR.n226 VDPWR.t357 44.3742
R1306 VDPWR.n446 VDPWR.t94 44.3742
R1307 VDPWR.n446 VDPWR.t405 44.3742
R1308 VDPWR.t78 VDPWR.n250 44.3742
R1309 VDPWR.n250 VDPWR.t51 44.3742
R1310 VDPWR.n420 VDPWR.t258 44.3742
R1311 VDPWR.n420 VDPWR.t256 44.3742
R1312 VDPWR.t554 VDPWR.n274 44.3742
R1313 VDPWR.n274 VDPWR.t274 44.3742
R1314 VDPWR.n394 VDPWR.t244 44.3742
R1315 VDPWR.n394 VDPWR.t355 44.3742
R1316 VDPWR.t123 VDPWR.n298 44.3742
R1317 VDPWR.n298 VDPWR.t514 44.3742
R1318 VDPWR.n368 VDPWR.t202 44.3742
R1319 VDPWR.n368 VDPWR.t412 44.3742
R1320 VDPWR.t420 VDPWR.n322 44.3742
R1321 VDPWR.n322 VDPWR.t435 44.3742
R1322 VDPWR.n334 VDPWR.t508 44.3742
R1323 VDPWR.n334 VDPWR.t351 44.3742
R1324 VDPWR.t449 VDPWR.n31 44.3742
R1325 VDPWR.n31 VDPWR.t423 44.3742
R1326 VDPWR.n101 VDPWR.t546 44.3742
R1327 VDPWR.n101 VDPWR.t277 44.3742
R1328 VDPWR.t417 VDPWR.n55 44.3742
R1329 VDPWR.n55 VDPWR.t432 44.3742
R1330 VDPWR.n67 VDPWR.t611 44.3742
R1331 VDPWR.n67 VDPWR.t609 44.3742
R1332 VDPWR.n181 VDPWR.n179 43.625
R1333 VDPWR.n175 VDPWR.n173 43.625
R1334 VDPWR.n10 VDPWR.n8 43.625
R1335 VDPWR.n4 VDPWR.n2 43.625
R1336 VDPWR.n507 VDPWR.n171 35.5442
R1337 VDPWR.n144 VDPWR.n0 35.5442
R1338 VDPWR.n496 VDPWR.n177 35.5275
R1339 VDPWR.n133 VDPWR.n6 35.5275
R1340 VDPWR.n530 VDPWR.n167 33.509
R1341 VDPWR.n1571 VDPWR.n1570 33.509
R1342 VDPWR.n520 VDPWR.n519 32.2656
R1343 VDPWR.n157 VDPWR.n156 32.2656
R1344 VDPWR.n579 VDPWR.n576 31.5192
R1345 VDPWR.n596 VDPWR.n593 31.5192
R1346 VDPWR.n613 VDPWR.n610 31.5192
R1347 VDPWR.n630 VDPWR.n627 31.5192
R1348 VDPWR.n647 VDPWR.n644 31.5192
R1349 VDPWR.n664 VDPWR.n661 31.5192
R1350 VDPWR.n681 VDPWR.n678 31.5192
R1351 VDPWR.n698 VDPWR.n695 31.5192
R1352 VDPWR.n188 VDPWR.t150 28.6437
R1353 VDPWR.n212 VDPWR.t527 28.6437
R1354 VDPWR.n236 VDPWR.t305 28.6437
R1355 VDPWR.n260 VDPWR.t74 28.6437
R1356 VDPWR.n284 VDPWR.t70 28.6437
R1357 VDPWR.n308 VDPWR.t254 28.6437
R1358 VDPWR.n17 VDPWR.t429 28.6437
R1359 VDPWR.n41 VDPWR.t137 28.6437
R1360 VDPWR.n467 VDPWR.n200 23.1255
R1361 VDPWR.n202 VDPWR.n200 23.1255
R1362 VDPWR.n474 VDPWR.n473 23.1255
R1363 VDPWR.n473 VDPWR.n472 23.1255
R1364 VDPWR.n441 VDPWR.n224 23.1255
R1365 VDPWR.n226 VDPWR.n224 23.1255
R1366 VDPWR.n448 VDPWR.n447 23.1255
R1367 VDPWR.n447 VDPWR.n446 23.1255
R1368 VDPWR.n415 VDPWR.n248 23.1255
R1369 VDPWR.n250 VDPWR.n248 23.1255
R1370 VDPWR.n422 VDPWR.n421 23.1255
R1371 VDPWR.n421 VDPWR.n420 23.1255
R1372 VDPWR.n389 VDPWR.n272 23.1255
R1373 VDPWR.n274 VDPWR.n272 23.1255
R1374 VDPWR.n396 VDPWR.n395 23.1255
R1375 VDPWR.n395 VDPWR.n394 23.1255
R1376 VDPWR.n363 VDPWR.n296 23.1255
R1377 VDPWR.n298 VDPWR.n296 23.1255
R1378 VDPWR.n370 VDPWR.n369 23.1255
R1379 VDPWR.n369 VDPWR.n368 23.1255
R1380 VDPWR.n329 VDPWR.n320 23.1255
R1381 VDPWR.n322 VDPWR.n320 23.1255
R1382 VDPWR.n336 VDPWR.n335 23.1255
R1383 VDPWR.n335 VDPWR.n334 23.1255
R1384 VDPWR.n96 VDPWR.n29 23.1255
R1385 VDPWR.n31 VDPWR.n29 23.1255
R1386 VDPWR.n103 VDPWR.n102 23.1255
R1387 VDPWR.n102 VDPWR.n101 23.1255
R1388 VDPWR.n62 VDPWR.n53 23.1255
R1389 VDPWR.n55 VDPWR.n53 23.1255
R1390 VDPWR.n69 VDPWR.n68 23.1255
R1391 VDPWR.n68 VDPWR.n67 23.1255
R1392 VDPWR.n495 VDPWR.t16 20.8338
R1393 VDPWR.n132 VDPWR.t0 20.8338
R1394 VDPWR.n506 VDPWR.t461 20.7429
R1395 VDPWR.n143 VDPWR.t474 20.7429
R1396 VDPWR.n1523 VDPWR.n1507 20.5561
R1397 VDPWR.n1540 VDPWR.n1523 20.5561
R1398 VDPWR.n1521 VDPWR.n1504 20.5561
R1399 VDPWR.n1540 VDPWR.n1521 20.5561
R1400 VDPWR.n1519 VDPWR.n1500 20.5561
R1401 VDPWR.n1540 VDPWR.n1519 20.5561
R1402 VDPWR.n1517 VDPWR.n1497 20.5561
R1403 VDPWR.n1540 VDPWR.n1517 20.5561
R1404 VDPWR.n1515 VDPWR.n1493 20.5561
R1405 VDPWR.n1540 VDPWR.n1515 20.5561
R1406 VDPWR.n1513 VDPWR.n1490 20.5561
R1407 VDPWR.n1540 VDPWR.n1513 20.5561
R1408 VDPWR.n1539 VDPWR.n1538 20.5561
R1409 VDPWR.n1540 VDPWR.n1539 20.5561
R1410 VDPWR.n1532 VDPWR.n1524 20.5561
R1411 VDPWR.n1540 VDPWR.n1524 20.5561
R1412 VDPWR.n1542 VDPWR.n1541 20.5561
R1413 VDPWR.n1541 VDPWR.n1540 20.5561
R1414 VDPWR.n1001 VDPWR.n1000 20.5561
R1415 VDPWR.n1004 VDPWR.n996 20.5561
R1416 VDPWR.n1005 VDPWR.n1004 20.5561
R1417 VDPWR.n1003 VDPWR.n994 20.5561
R1418 VDPWR.n1019 VDPWR.n1018 20.5561
R1419 VDPWR.n1022 VDPWR.n992 20.5561
R1420 VDPWR.n1023 VDPWR.n1022 20.5561
R1421 VDPWR.n1021 VDPWR.n990 20.5561
R1422 VDPWR.n1037 VDPWR.n1036 20.5561
R1423 VDPWR.n1040 VDPWR.n988 20.5561
R1424 VDPWR.n1041 VDPWR.n1040 20.5561
R1425 VDPWR.n1039 VDPWR.n986 20.5561
R1426 VDPWR.n1055 VDPWR.n1054 20.5561
R1427 VDPWR.n1058 VDPWR.n984 20.5561
R1428 VDPWR.n1059 VDPWR.n1058 20.5561
R1429 VDPWR.n1057 VDPWR.n982 20.5561
R1430 VDPWR.n1073 VDPWR.n1072 20.5561
R1431 VDPWR.n1076 VDPWR.n980 20.5561
R1432 VDPWR.n1077 VDPWR.n1076 20.5561
R1433 VDPWR.n1075 VDPWR.n978 20.5561
R1434 VDPWR.n1091 VDPWR.n1090 20.5561
R1435 VDPWR.n1094 VDPWR.n976 20.5561
R1436 VDPWR.n1095 VDPWR.n1094 20.5561
R1437 VDPWR.n1093 VDPWR.n974 20.5561
R1438 VDPWR.n1109 VDPWR.n1108 20.5561
R1439 VDPWR.n1112 VDPWR.n972 20.5561
R1440 VDPWR.n1113 VDPWR.n1112 20.5561
R1441 VDPWR.n1111 VDPWR.n970 20.5561
R1442 VDPWR.n1127 VDPWR.n1126 20.5561
R1443 VDPWR.n1130 VDPWR.n968 20.5561
R1444 VDPWR.n1131 VDPWR.n1130 20.5561
R1445 VDPWR.n1129 VDPWR.n966 20.5561
R1446 VDPWR.n857 VDPWR.n798 20.5561
R1447 VDPWR.n863 VDPWR.n857 20.5561
R1448 VDPWR.n855 VDPWR.n795 20.5561
R1449 VDPWR.n863 VDPWR.n855 20.5561
R1450 VDPWR.n853 VDPWR.n791 20.5561
R1451 VDPWR.n863 VDPWR.n853 20.5561
R1452 VDPWR.n851 VDPWR.n788 20.5561
R1453 VDPWR.n863 VDPWR.n851 20.5561
R1454 VDPWR.n849 VDPWR.n784 20.5561
R1455 VDPWR.n863 VDPWR.n849 20.5561
R1456 VDPWR.n847 VDPWR.n781 20.5561
R1457 VDPWR.n863 VDPWR.n847 20.5561
R1458 VDPWR.n845 VDPWR.n777 20.5561
R1459 VDPWR.n863 VDPWR.n845 20.5561
R1460 VDPWR.n843 VDPWR.n774 20.5561
R1461 VDPWR.n863 VDPWR.n843 20.5561
R1462 VDPWR.n841 VDPWR.n770 20.5561
R1463 VDPWR.n863 VDPWR.n841 20.5561
R1464 VDPWR.n839 VDPWR.n767 20.5561
R1465 VDPWR.n863 VDPWR.n839 20.5561
R1466 VDPWR.n837 VDPWR.n763 20.5561
R1467 VDPWR.n863 VDPWR.n837 20.5561
R1468 VDPWR.n835 VDPWR.n760 20.5561
R1469 VDPWR.n863 VDPWR.n835 20.5561
R1470 VDPWR.n833 VDPWR.n756 20.5561
R1471 VDPWR.n863 VDPWR.n833 20.5561
R1472 VDPWR.n831 VDPWR.n753 20.5561
R1473 VDPWR.n863 VDPWR.n831 20.5561
R1474 VDPWR.n829 VDPWR.n749 20.5561
R1475 VDPWR.n863 VDPWR.n829 20.5561
R1476 VDPWR.n827 VDPWR.n746 20.5561
R1477 VDPWR.n863 VDPWR.n827 20.5561
R1478 VDPWR.n825 VDPWR.n742 20.5561
R1479 VDPWR.n863 VDPWR.n825 20.5561
R1480 VDPWR.n823 VDPWR.n739 20.5561
R1481 VDPWR.n863 VDPWR.n823 20.5561
R1482 VDPWR.n821 VDPWR.n735 20.5561
R1483 VDPWR.n863 VDPWR.n821 20.5561
R1484 VDPWR.n819 VDPWR.n732 20.5561
R1485 VDPWR.n863 VDPWR.n819 20.5561
R1486 VDPWR.n817 VDPWR.n728 20.5561
R1487 VDPWR.n863 VDPWR.n817 20.5561
R1488 VDPWR.n815 VDPWR.n725 20.5561
R1489 VDPWR.n863 VDPWR.n815 20.5561
R1490 VDPWR.n813 VDPWR.n721 20.5561
R1491 VDPWR.n863 VDPWR.n813 20.5561
R1492 VDPWR.n811 VDPWR.n718 20.5561
R1493 VDPWR.n863 VDPWR.n811 20.5561
R1494 VDPWR.n809 VDPWR.n714 20.5561
R1495 VDPWR.n863 VDPWR.n809 20.5561
R1496 VDPWR.n807 VDPWR.n711 20.5561
R1497 VDPWR.n863 VDPWR.n807 20.5561
R1498 VDPWR.n862 VDPWR.n802 20.5561
R1499 VDPWR.n863 VDPWR.n862 20.5561
R1500 VDPWR.n859 VDPWR.n805 20.5561
R1501 VDPWR.n863 VDPWR.n859 20.5561
R1502 VDPWR.n865 VDPWR.n864 20.5561
R1503 VDPWR.n864 VDPWR.n863 20.5561
R1504 VDPWR.n517 VDPWR.n514 20.5561
R1505 VDPWR.n518 VDPWR.n517 20.5561
R1506 VDPWR.n494 VDPWR.n493 20.5561
R1507 VDPWR.n495 VDPWR.n494 20.5561
R1508 VDPWR.n182 VDPWR.n181 20.5561
R1509 VDPWR.n495 VDPWR.n182 20.5561
R1510 VDPWR.n505 VDPWR.n504 20.5561
R1511 VDPWR.n506 VDPWR.n505 20.5561
R1512 VDPWR.n176 VDPWR.n175 20.5561
R1513 VDPWR.n506 VDPWR.n176 20.5561
R1514 VDPWR.n192 VDPWR.n190 20.5561
R1515 VDPWR.n190 VDPWR.n188 20.5561
R1516 VDPWR.n191 VDPWR.n189 20.5561
R1517 VDPWR.n189 VDPWR.n188 20.5561
R1518 VDPWR.n186 VDPWR.n185 20.5561
R1519 VDPWR.n188 VDPWR.n186 20.5561
R1520 VDPWR.n187 VDPWR.n183 20.5561
R1521 VDPWR.n188 VDPWR.n187 20.5561
R1522 VDPWR.n216 VDPWR.n214 20.5561
R1523 VDPWR.n214 VDPWR.n212 20.5561
R1524 VDPWR.n215 VDPWR.n213 20.5561
R1525 VDPWR.n213 VDPWR.n212 20.5561
R1526 VDPWR.n210 VDPWR.n209 20.5561
R1527 VDPWR.n212 VDPWR.n210 20.5561
R1528 VDPWR.n211 VDPWR.n207 20.5561
R1529 VDPWR.n212 VDPWR.n211 20.5561
R1530 VDPWR.n240 VDPWR.n238 20.5561
R1531 VDPWR.n238 VDPWR.n236 20.5561
R1532 VDPWR.n239 VDPWR.n237 20.5561
R1533 VDPWR.n237 VDPWR.n236 20.5561
R1534 VDPWR.n234 VDPWR.n233 20.5561
R1535 VDPWR.n236 VDPWR.n234 20.5561
R1536 VDPWR.n235 VDPWR.n231 20.5561
R1537 VDPWR.n236 VDPWR.n235 20.5561
R1538 VDPWR.n264 VDPWR.n262 20.5561
R1539 VDPWR.n262 VDPWR.n260 20.5561
R1540 VDPWR.n263 VDPWR.n261 20.5561
R1541 VDPWR.n261 VDPWR.n260 20.5561
R1542 VDPWR.n258 VDPWR.n257 20.5561
R1543 VDPWR.n260 VDPWR.n258 20.5561
R1544 VDPWR.n259 VDPWR.n255 20.5561
R1545 VDPWR.n260 VDPWR.n259 20.5561
R1546 VDPWR.n288 VDPWR.n286 20.5561
R1547 VDPWR.n286 VDPWR.n284 20.5561
R1548 VDPWR.n287 VDPWR.n285 20.5561
R1549 VDPWR.n285 VDPWR.n284 20.5561
R1550 VDPWR.n282 VDPWR.n281 20.5561
R1551 VDPWR.n284 VDPWR.n282 20.5561
R1552 VDPWR.n283 VDPWR.n279 20.5561
R1553 VDPWR.n284 VDPWR.n283 20.5561
R1554 VDPWR.n312 VDPWR.n310 20.5561
R1555 VDPWR.n310 VDPWR.n308 20.5561
R1556 VDPWR.n311 VDPWR.n309 20.5561
R1557 VDPWR.n309 VDPWR.n308 20.5561
R1558 VDPWR.n306 VDPWR.n305 20.5561
R1559 VDPWR.n308 VDPWR.n306 20.5561
R1560 VDPWR.n307 VDPWR.n303 20.5561
R1561 VDPWR.n308 VDPWR.n307 20.5561
R1562 VDPWR.n528 VDPWR.n527 20.5561
R1563 VDPWR.n529 VDPWR.n528 20.5561
R1564 VDPWR.n154 VDPWR.n151 20.5561
R1565 VDPWR.n155 VDPWR.n154 20.5561
R1566 VDPWR.n131 VDPWR.n130 20.5561
R1567 VDPWR.n132 VDPWR.n131 20.5561
R1568 VDPWR.n11 VDPWR.n10 20.5561
R1569 VDPWR.n132 VDPWR.n11 20.5561
R1570 VDPWR.n142 VDPWR.n141 20.5561
R1571 VDPWR.n143 VDPWR.n142 20.5561
R1572 VDPWR.n5 VDPWR.n4 20.5561
R1573 VDPWR.n143 VDPWR.n5 20.5561
R1574 VDPWR.n21 VDPWR.n19 20.5561
R1575 VDPWR.n19 VDPWR.n17 20.5561
R1576 VDPWR.n20 VDPWR.n18 20.5561
R1577 VDPWR.n18 VDPWR.n17 20.5561
R1578 VDPWR.n15 VDPWR.n14 20.5561
R1579 VDPWR.n17 VDPWR.n15 20.5561
R1580 VDPWR.n16 VDPWR.n12 20.5561
R1581 VDPWR.n17 VDPWR.n16 20.5561
R1582 VDPWR.n40 VDPWR.n36 20.5561
R1583 VDPWR.n41 VDPWR.n40 20.5561
R1584 VDPWR.n39 VDPWR.n38 20.5561
R1585 VDPWR.n41 VDPWR.n39 20.5561
R1586 VDPWR.n45 VDPWR.n43 20.5561
R1587 VDPWR.n43 VDPWR.n41 20.5561
R1588 VDPWR.n44 VDPWR.n42 20.5561
R1589 VDPWR.n42 VDPWR.n41 20.5561
R1590 VDPWR.n1574 VDPWR.n1573 20.5561
R1591 VDPWR.n1573 VDPWR.n1572 20.5561
R1592 VDPWR.n1562 VDPWR.n1561 19.3338
R1593 VDPWR.n1561 VDPWR.n1560 19.3338
R1594 VDPWR.n1560 VDPWR.n1495 19.3338
R1595 VDPWR.n1555 VDPWR.n1495 19.3338
R1596 VDPWR.n1555 VDPWR.n1554 19.3338
R1597 VDPWR.n1554 VDPWR.n1553 19.3338
R1598 VDPWR.n1553 VDPWR.n1502 19.3338
R1599 VDPWR.n1548 VDPWR.n1502 19.3338
R1600 VDPWR.n1548 VDPWR.n1547 19.3338
R1601 VDPWR.n1547 VDPWR.n1546 19.3338
R1602 VDPWR.n1546 VDPWR.n1509 19.3338
R1603 VDPWR.n1530 VDPWR.n1509 19.3338
R1604 VDPWR.n1537 VDPWR.n1530 19.3338
R1605 VDPWR.n1537 VDPWR.n1536 19.3338
R1606 VDPWR.n963 VDPWR.n962 19.3338
R1607 VDPWR.n962 VDPWR.n961 19.3338
R1608 VDPWR.n961 VDPWR.n716 19.3338
R1609 VDPWR.n956 VDPWR.n716 19.3338
R1610 VDPWR.n956 VDPWR.n955 19.3338
R1611 VDPWR.n955 VDPWR.n954 19.3338
R1612 VDPWR.n954 VDPWR.n723 19.3338
R1613 VDPWR.n949 VDPWR.n723 19.3338
R1614 VDPWR.n949 VDPWR.n948 19.3338
R1615 VDPWR.n948 VDPWR.n947 19.3338
R1616 VDPWR.n947 VDPWR.n730 19.3338
R1617 VDPWR.n942 VDPWR.n730 19.3338
R1618 VDPWR.n942 VDPWR.n941 19.3338
R1619 VDPWR.n941 VDPWR.n940 19.3338
R1620 VDPWR.n940 VDPWR.n737 19.3338
R1621 VDPWR.n935 VDPWR.n737 19.3338
R1622 VDPWR.n935 VDPWR.n934 19.3338
R1623 VDPWR.n934 VDPWR.n933 19.3338
R1624 VDPWR.n933 VDPWR.n744 19.3338
R1625 VDPWR.n928 VDPWR.n744 19.3338
R1626 VDPWR.n928 VDPWR.n927 19.3338
R1627 VDPWR.n927 VDPWR.n926 19.3338
R1628 VDPWR.n926 VDPWR.n751 19.3338
R1629 VDPWR.n921 VDPWR.n751 19.3338
R1630 VDPWR.n921 VDPWR.n920 19.3338
R1631 VDPWR.n920 VDPWR.n919 19.3338
R1632 VDPWR.n919 VDPWR.n758 19.3338
R1633 VDPWR.n914 VDPWR.n758 19.3338
R1634 VDPWR.n914 VDPWR.n913 19.3338
R1635 VDPWR.n913 VDPWR.n912 19.3338
R1636 VDPWR.n912 VDPWR.n765 19.3338
R1637 VDPWR.n907 VDPWR.n765 19.3338
R1638 VDPWR.n907 VDPWR.n906 19.3338
R1639 VDPWR.n906 VDPWR.n905 19.3338
R1640 VDPWR.n905 VDPWR.n772 19.3338
R1641 VDPWR.n900 VDPWR.n772 19.3338
R1642 VDPWR.n900 VDPWR.n899 19.3338
R1643 VDPWR.n899 VDPWR.n898 19.3338
R1644 VDPWR.n898 VDPWR.n779 19.3338
R1645 VDPWR.n893 VDPWR.n779 19.3338
R1646 VDPWR.n893 VDPWR.n892 19.3338
R1647 VDPWR.n892 VDPWR.n891 19.3338
R1648 VDPWR.n891 VDPWR.n786 19.3338
R1649 VDPWR.n886 VDPWR.n786 19.3338
R1650 VDPWR.n886 VDPWR.n885 19.3338
R1651 VDPWR.n885 VDPWR.n884 19.3338
R1652 VDPWR.n884 VDPWR.n793 19.3338
R1653 VDPWR.n879 VDPWR.n793 19.3338
R1654 VDPWR.n879 VDPWR.n878 19.3338
R1655 VDPWR.n878 VDPWR.n877 19.3338
R1656 VDPWR.n877 VDPWR.n800 19.3338
R1657 VDPWR.n872 VDPWR.n800 19.3338
R1658 VDPWR.n872 VDPWR.n871 19.3338
R1659 VDPWR.n871 VDPWR.n870 19.3338
R1660 VDPWR.n702 VDPWR.n700 18.5005
R1661 VDPWR.n706 VDPWR.n700 18.5005
R1662 VDPWR.n685 VDPWR.n683 18.5005
R1663 VDPWR.n689 VDPWR.n683 18.5005
R1664 VDPWR.n668 VDPWR.n666 18.5005
R1665 VDPWR.n672 VDPWR.n666 18.5005
R1666 VDPWR.n651 VDPWR.n649 18.5005
R1667 VDPWR.n655 VDPWR.n649 18.5005
R1668 VDPWR.n634 VDPWR.n632 18.5005
R1669 VDPWR.n638 VDPWR.n632 18.5005
R1670 VDPWR.n617 VDPWR.n615 18.5005
R1671 VDPWR.n621 VDPWR.n615 18.5005
R1672 VDPWR.n600 VDPWR.n598 18.5005
R1673 VDPWR.n604 VDPWR.n598 18.5005
R1674 VDPWR.n583 VDPWR.n581 18.5005
R1675 VDPWR.n587 VDPWR.n581 18.5005
R1676 VDPWR.n589 VDPWR.n588 18.5005
R1677 VDPWR.n588 VDPWR.n587 18.5005
R1678 VDPWR.n606 VDPWR.n605 18.5005
R1679 VDPWR.n605 VDPWR.n604 18.5005
R1680 VDPWR.n623 VDPWR.n622 18.5005
R1681 VDPWR.n622 VDPWR.n621 18.5005
R1682 VDPWR.n640 VDPWR.n639 18.5005
R1683 VDPWR.n639 VDPWR.n638 18.5005
R1684 VDPWR.n657 VDPWR.n656 18.5005
R1685 VDPWR.n656 VDPWR.n655 18.5005
R1686 VDPWR.n674 VDPWR.n673 18.5005
R1687 VDPWR.n673 VDPWR.n672 18.5005
R1688 VDPWR.n691 VDPWR.n690 18.5005
R1689 VDPWR.n690 VDPWR.n689 18.5005
R1690 VDPWR.n708 VDPWR.n707 18.5005
R1691 VDPWR.n707 VDPWR.n706 18.5005
R1692 VDPWR.n469 VDPWR.n468 18.5005
R1693 VDPWR.n470 VDPWR.n469 18.5005
R1694 VDPWR.n204 VDPWR.n203 18.5005
R1695 VDPWR.n198 VDPWR.n197 18.5005
R1696 VDPWR.n471 VDPWR.n198 18.5005
R1697 VDPWR.n199 VDPWR.n193 18.5005
R1698 VDPWR.n443 VDPWR.n442 18.5005
R1699 VDPWR.n444 VDPWR.n443 18.5005
R1700 VDPWR.n228 VDPWR.n227 18.5005
R1701 VDPWR.n222 VDPWR.n221 18.5005
R1702 VDPWR.n445 VDPWR.n222 18.5005
R1703 VDPWR.n223 VDPWR.n217 18.5005
R1704 VDPWR.n417 VDPWR.n416 18.5005
R1705 VDPWR.n418 VDPWR.n417 18.5005
R1706 VDPWR.n252 VDPWR.n251 18.5005
R1707 VDPWR.n246 VDPWR.n245 18.5005
R1708 VDPWR.n419 VDPWR.n246 18.5005
R1709 VDPWR.n247 VDPWR.n241 18.5005
R1710 VDPWR.n391 VDPWR.n390 18.5005
R1711 VDPWR.n392 VDPWR.n391 18.5005
R1712 VDPWR.n276 VDPWR.n275 18.5005
R1713 VDPWR.n270 VDPWR.n269 18.5005
R1714 VDPWR.n393 VDPWR.n270 18.5005
R1715 VDPWR.n271 VDPWR.n265 18.5005
R1716 VDPWR.n365 VDPWR.n364 18.5005
R1717 VDPWR.n366 VDPWR.n365 18.5005
R1718 VDPWR.n300 VDPWR.n299 18.5005
R1719 VDPWR.n294 VDPWR.n293 18.5005
R1720 VDPWR.n367 VDPWR.n294 18.5005
R1721 VDPWR.n295 VDPWR.n289 18.5005
R1722 VDPWR.n331 VDPWR.n330 18.5005
R1723 VDPWR.n332 VDPWR.n331 18.5005
R1724 VDPWR.n324 VDPWR.n323 18.5005
R1725 VDPWR.n318 VDPWR.n317 18.5005
R1726 VDPWR.n333 VDPWR.n318 18.5005
R1727 VDPWR.n319 VDPWR.n313 18.5005
R1728 VDPWR.n532 VDPWR.n531 18.5005
R1729 VDPWR.n98 VDPWR.n97 18.5005
R1730 VDPWR.n99 VDPWR.n98 18.5005
R1731 VDPWR.n33 VDPWR.n32 18.5005
R1732 VDPWR.n27 VDPWR.n26 18.5005
R1733 VDPWR.n100 VDPWR.n27 18.5005
R1734 VDPWR.n28 VDPWR.n22 18.5005
R1735 VDPWR.n64 VDPWR.n63 18.5005
R1736 VDPWR.n65 VDPWR.n64 18.5005
R1737 VDPWR.n57 VDPWR.n56 18.5005
R1738 VDPWR.n51 VDPWR.n50 18.5005
R1739 VDPWR.n66 VDPWR.n51 18.5005
R1740 VDPWR.n52 VDPWR.n46 18.5005
R1741 VDPWR.n164 VDPWR.n163 18.5005
R1742 VDPWR.n1194 VDPWR.n1193 16.8187
R1743 VDPWR.n1196 VDPWR.n1195 16.8187
R1744 VDPWR.n1190 VDPWR.n1183 16.8187
R1745 VDPWR.n1197 VDPWR.n1190 16.8187
R1746 VDPWR.n1210 VDPWR.n1208 16.8187
R1747 VDPWR.n1211 VDPWR.n1178 16.8187
R1748 VDPWR.n1212 VDPWR.n1211 16.8187
R1749 VDPWR.n1226 VDPWR.n1224 16.8187
R1750 VDPWR.n1227 VDPWR.n1173 16.8187
R1751 VDPWR.n1228 VDPWR.n1227 16.8187
R1752 VDPWR.n1242 VDPWR.n1240 16.8187
R1753 VDPWR.n1243 VDPWR.n1168 16.8187
R1754 VDPWR.n1244 VDPWR.n1243 16.8187
R1755 VDPWR.n1258 VDPWR.n1256 16.8187
R1756 VDPWR.n1259 VDPWR.n1163 16.8187
R1757 VDPWR.n1260 VDPWR.n1259 16.8187
R1758 VDPWR.n1274 VDPWR.n1272 16.8187
R1759 VDPWR.n1275 VDPWR.n1158 16.8187
R1760 VDPWR.n1276 VDPWR.n1275 16.8187
R1761 VDPWR.n1290 VDPWR.n1288 16.8187
R1762 VDPWR.n1291 VDPWR.n1153 16.8187
R1763 VDPWR.n1292 VDPWR.n1291 16.8187
R1764 VDPWR.n1306 VDPWR.n1304 16.8187
R1765 VDPWR.n1307 VDPWR.n1148 16.8187
R1766 VDPWR.n1308 VDPWR.n1307 16.8187
R1767 VDPWR.n1322 VDPWR.n1320 16.8187
R1768 VDPWR.n1323 VDPWR.n1143 16.8187
R1769 VDPWR.n1324 VDPWR.n1323 16.8187
R1770 VDPWR.n590 VDPWR.n575 16.8187
R1771 VDPWR.n578 VDPWR.n575 16.8187
R1772 VDPWR.n607 VDPWR.n570 16.8187
R1773 VDPWR.n595 VDPWR.n570 16.8187
R1774 VDPWR.n624 VDPWR.n565 16.8187
R1775 VDPWR.n612 VDPWR.n565 16.8187
R1776 VDPWR.n641 VDPWR.n560 16.8187
R1777 VDPWR.n629 VDPWR.n560 16.8187
R1778 VDPWR.n658 VDPWR.n555 16.8187
R1779 VDPWR.n646 VDPWR.n555 16.8187
R1780 VDPWR.n675 VDPWR.n550 16.8187
R1781 VDPWR.n663 VDPWR.n550 16.8187
R1782 VDPWR.n692 VDPWR.n545 16.8187
R1783 VDPWR.n680 VDPWR.n545 16.8187
R1784 VDPWR.n709 VDPWR.n540 16.8187
R1785 VDPWR.n697 VDPWR.n540 16.8187
R1786 VDPWR.n1480 VDPWR.n1335 16.8187
R1787 VDPWR.n1481 VDPWR.n1480 16.8187
R1788 VDPWR.n1478 VDPWR.n1340 16.8187
R1789 VDPWR.n1479 VDPWR.n1478 16.8187
R1790 VDPWR.n1476 VDPWR.n1475 16.8187
R1791 VDPWR.n1477 VDPWR.n1476 16.8187
R1792 VDPWR.n1454 VDPWR.n1347 16.8187
R1793 VDPWR.n1455 VDPWR.n1454 16.8187
R1794 VDPWR.n1456 VDPWR.n1351 16.8187
R1795 VDPWR.n1457 VDPWR.n1456 16.8187
R1796 VDPWR.n1450 VDPWR.n1356 16.8187
R1797 VDPWR.n1451 VDPWR.n1450 16.8187
R1798 VDPWR.n1448 VDPWR.n1447 16.8187
R1799 VDPWR.n1449 VDPWR.n1448 16.8187
R1800 VDPWR.n1426 VDPWR.n1363 16.8187
R1801 VDPWR.n1427 VDPWR.n1426 16.8187
R1802 VDPWR.n1428 VDPWR.n1367 16.8187
R1803 VDPWR.n1429 VDPWR.n1428 16.8187
R1804 VDPWR.n1422 VDPWR.n1372 16.8187
R1805 VDPWR.n1423 VDPWR.n1422 16.8187
R1806 VDPWR.n1420 VDPWR.n1419 16.8187
R1807 VDPWR.n1421 VDPWR.n1420 16.8187
R1808 VDPWR.n1400 VDPWR.n1379 16.8187
R1809 VDPWR.n1401 VDPWR.n1400 16.8187
R1810 VDPWR.n1397 VDPWR.n1396 16.8187
R1811 VDPWR.n1390 VDPWR.n1383 16.8187
R1812 VDPWR.n1402 VDPWR.n1390 16.8187
R1813 VDPWR.n1395 VDPWR.n1394 16.8187
R1814 VDPWR.n589 VDPWR.n576 14.3397
R1815 VDPWR.n606 VDPWR.n593 14.3397
R1816 VDPWR.n623 VDPWR.n610 14.3397
R1817 VDPWR.n640 VDPWR.n627 14.3397
R1818 VDPWR.n657 VDPWR.n644 14.3397
R1819 VDPWR.n674 VDPWR.n661 14.3397
R1820 VDPWR.n691 VDPWR.n678 14.3397
R1821 VDPWR.n708 VDPWR.n695 14.3397
R1822 VDPWR.n704 VDPWR.n702 13.8537
R1823 VDPWR.n702 VDPWR.n695 13.8537
R1824 VDPWR.n687 VDPWR.n685 13.8537
R1825 VDPWR.n685 VDPWR.n678 13.8537
R1826 VDPWR.n670 VDPWR.n668 13.8537
R1827 VDPWR.n668 VDPWR.n661 13.8537
R1828 VDPWR.n653 VDPWR.n651 13.8537
R1829 VDPWR.n651 VDPWR.n644 13.8537
R1830 VDPWR.n636 VDPWR.n634 13.8537
R1831 VDPWR.n634 VDPWR.n627 13.8537
R1832 VDPWR.n619 VDPWR.n617 13.8537
R1833 VDPWR.n617 VDPWR.n610 13.8537
R1834 VDPWR.n602 VDPWR.n600 13.8537
R1835 VDPWR.n600 VDPWR.n593 13.8537
R1836 VDPWR.n585 VDPWR.n583 13.8537
R1837 VDPWR.n583 VDPWR.n576 13.8537
R1838 VDPWR.n703 VDPWR.n699 13.2148
R1839 VDPWR.n686 VDPWR.n682 13.2148
R1840 VDPWR.n669 VDPWR.n665 13.2148
R1841 VDPWR.n652 VDPWR.n648 13.2148
R1842 VDPWR.n635 VDPWR.n631 13.2148
R1843 VDPWR.n618 VDPWR.n614 13.2148
R1844 VDPWR.n601 VDPWR.n597 13.2148
R1845 VDPWR.n584 VDPWR.n580 13.2148
R1846 VDPWR.n1200 VDPWR.n1199 11.563
R1847 VDPWR.n1199 VDPWR.n1198 11.563
R1848 VDPWR.n1213 VDPWR.n1209 11.563
R1849 VDPWR.n1229 VDPWR.n1225 11.563
R1850 VDPWR.n1245 VDPWR.n1241 11.563
R1851 VDPWR.n1261 VDPWR.n1257 11.563
R1852 VDPWR.n1277 VDPWR.n1273 11.563
R1853 VDPWR.n1293 VDPWR.n1289 11.563
R1854 VDPWR.n1309 VDPWR.n1305 11.563
R1855 VDPWR.n1325 VDPWR.n1321 11.563
R1856 VDPWR.n1482 VDPWR.n1341 11.563
R1857 VDPWR.n1452 VDPWR.n1342 11.563
R1858 VDPWR.n1458 VDPWR.n1357 11.563
R1859 VDPWR.n1424 VDPWR.n1358 11.563
R1860 VDPWR.n1430 VDPWR.n1373 11.563
R1861 VDPWR.n1398 VDPWR.n1374 11.563
R1862 VDPWR.n1405 VDPWR.n1404 11.563
R1863 VDPWR.n1404 VDPWR.n1403 11.563
R1864 VDPWR.n1215 VDPWR.n1209 10.2708
R1865 VDPWR.n1231 VDPWR.n1225 10.2708
R1866 VDPWR.n1247 VDPWR.n1241 10.2708
R1867 VDPWR.n1263 VDPWR.n1257 10.2708
R1868 VDPWR.n1279 VDPWR.n1273 10.2708
R1869 VDPWR.n1295 VDPWR.n1289 10.2708
R1870 VDPWR.n1311 VDPWR.n1305 10.2708
R1871 VDPWR.n1327 VDPWR.n1321 10.2708
R1872 VDPWR.n1484 VDPWR.n1341 10.2708
R1873 VDPWR.n1348 VDPWR.n1342 10.2708
R1874 VDPWR.n1460 VDPWR.n1357 10.2708
R1875 VDPWR.n1364 VDPWR.n1358 10.2708
R1876 VDPWR.n1432 VDPWR.n1373 10.2708
R1877 VDPWR.n1380 VDPWR.n1374 10.2708
R1878 VDPWR.n1386 VDPWR.t376 9.52217
R1879 VDPWR.n1386 VDPWR.t518 9.52217
R1880 VDPWR.n1385 VDPWR.t147 9.52217
R1881 VDPWR.n1385 VDPWR.t11 9.52217
R1882 VDPWR.n1384 VDPWR.t9 9.52217
R1883 VDPWR.n1384 VDPWR.t34 9.52217
R1884 VDPWR.n1382 VDPWR.t316 9.52217
R1885 VDPWR.n1382 VDPWR.t142 9.52217
R1886 VDPWR.n1381 VDPWR.t591 9.52217
R1887 VDPWR.n1381 VDPWR.t314 9.52217
R1888 VDPWR.n1413 VDPWR.t308 9.52217
R1889 VDPWR.n1413 VDPWR.t310 9.52217
R1890 VDPWR.n1414 VDPWR.t497 9.52217
R1891 VDPWR.n1414 VDPWR.t312 9.52217
R1892 VDPWR.n1375 VDPWR.t559 9.52217
R1893 VDPWR.n1375 VDPWR.t557 9.52217
R1894 VDPWR.n1370 VDPWR.t261 9.52217
R1895 VDPWR.n1370 VDPWR.t561 9.52217
R1896 VDPWR.n1369 VDPWR.t545 9.52217
R1897 VDPWR.n1369 VDPWR.t323 9.52217
R1898 VDPWR.n1368 VDPWR.t387 9.52217
R1899 VDPWR.n1368 VDPWR.t144 9.52217
R1900 VDPWR.n1366 VDPWR.t488 9.52217
R1901 VDPWR.n1366 VDPWR.t464 9.52217
R1902 VDPWR.n1365 VDPWR.t237 9.52217
R1903 VDPWR.n1365 VDPWR.t209 9.52217
R1904 VDPWR.n1441 VDPWR.t364 9.52217
R1905 VDPWR.n1441 VDPWR.t368 9.52217
R1906 VDPWR.n1442 VDPWR.t366 9.52217
R1907 VDPWR.n1442 VDPWR.t472 9.52217
R1908 VDPWR.n1359 VDPWR.t321 9.52217
R1909 VDPWR.n1359 VDPWR.t140 9.52217
R1910 VDPWR.n1354 VDPWR.t374 9.52217
R1911 VDPWR.n1354 VDPWR.t543 9.52217
R1912 VDPWR.n1353 VDPWR.t495 9.52217
R1913 VDPWR.n1353 VDPWR.t616 9.52217
R1914 VDPWR.n1352 VDPWR.t220 9.52217
R1915 VDPWR.n1352 VDPWR.t520 9.52217
R1916 VDPWR.n1350 VDPWR.t129 9.52217
R1917 VDPWR.n1350 VDPWR.t271 9.52217
R1918 VDPWR.n1349 VDPWR.t501 9.52217
R1919 VDPWR.n1349 VDPWR.t73 9.52217
R1920 VDPWR.n1469 VDPWR.t179 9.52217
R1921 VDPWR.n1469 VDPWR.t470 9.52217
R1922 VDPWR.n1470 VDPWR.t468 9.52217
R1923 VDPWR.n1470 VDPWR.t181 9.52217
R1924 VDPWR.n1343 VDPWR.t253 9.52217
R1925 VDPWR.n1343 VDPWR.t91 9.52217
R1926 VDPWR.n1338 VDPWR.t249 9.52217
R1927 VDPWR.n1338 VDPWR.t251 9.52217
R1928 VDPWR.n1337 VDPWR.t36 9.52217
R1929 VDPWR.n1337 VDPWR.t44 9.52217
R1930 VDPWR.n1336 VDPWR.t46 9.52217
R1931 VDPWR.n1336 VDPWR.t404 9.52217
R1932 VDPWR.n1191 VDPWR.t507 9.52217
R1933 VDPWR.n1191 VDPWR.t466 9.52217
R1934 VDPWR.n1186 VDPWR.t393 9.52217
R1935 VDPWR.n1186 VDPWR.t350 9.52217
R1936 VDPWR.n1185 VDPWR.t571 9.52217
R1937 VDPWR.n1185 VDPWR.t269 9.52217
R1938 VDPWR.n1184 VDPWR.t333 9.52217
R1939 VDPWR.n1184 VDPWR.t331 9.52217
R1940 VDPWR.n1205 VDPWR.t551 9.52217
R1941 VDPWR.n1205 VDPWR.t177 9.52217
R1942 VDPWR.n1181 VDPWR.t175 9.52217
R1943 VDPWR.n1181 VDPWR.t190 9.52217
R1944 VDPWR.n1180 VDPWR.t67 9.52217
R1945 VDPWR.n1180 VDPWR.t65 9.52217
R1946 VDPWR.n1179 VDPWR.t541 9.52217
R1947 VDPWR.n1179 VDPWR.t587 9.52217
R1948 VDPWR.n1221 VDPWR.t288 9.52217
R1949 VDPWR.n1221 VDPWR.t297 9.52217
R1950 VDPWR.n1176 VDPWR.t218 9.52217
R1951 VDPWR.n1176 VDPWR.t207 9.52217
R1952 VDPWR.n1175 VDPWR.t399 9.52217
R1953 VDPWR.n1175 VDPWR.t524 9.52217
R1954 VDPWR.n1174 VDPWR.t522 9.52217
R1955 VDPWR.n1174 VDPWR.t31 9.52217
R1956 VDPWR.n1237 VDPWR.t411 9.52217
R1957 VDPWR.n1237 VDPWR.t48 9.52217
R1958 VDPWR.n1171 VDPWR.t93 9.52217
R1959 VDPWR.n1171 VDPWR.t578 9.52217
R1960 VDPWR.n1170 VDPWR.t604 9.52217
R1961 VDPWR.n1170 VDPWR.t60 9.52217
R1962 VDPWR.n1169 VDPWR.t391 9.52217
R1963 VDPWR.n1169 VDPWR.t163 9.52217
R1964 VDPWR.n1253 VDPWR.t183 9.52217
R1965 VDPWR.n1253 VDPWR.t481 9.52217
R1966 VDPWR.n1166 VDPWR.t282 9.52217
R1967 VDPWR.n1166 VDPWR.t280 9.52217
R1968 VDPWR.n1165 VDPWR.t87 9.52217
R1969 VDPWR.n1165 VDPWR.t499 9.52217
R1970 VDPWR.n1164 VDPWR.t247 9.52217
R1971 VDPWR.n1164 VDPWR.t168 9.52217
R1972 VDPWR.n1269 VDPWR.t460 9.52217
R1973 VDPWR.n1269 VDPWR.t454 9.52217
R1974 VDPWR.n1161 VDPWR.t456 9.52217
R1975 VDPWR.n1161 VDPWR.t458 9.52217
R1976 VDPWR.n1160 VDPWR.t329 9.52217
R1977 VDPWR.n1160 VDPWR.t362 9.52217
R1978 VDPWR.n1159 VDPWR.t378 9.52217
R1979 VDPWR.n1159 VDPWR.t360 9.52217
R1980 VDPWR.n1285 VDPWR.t113 9.52217
R1981 VDPWR.n1285 VDPWR.t409 9.52217
R1982 VDPWR.n1156 VDPWR.t372 9.52217
R1983 VDPWR.n1156 VDPWR.t370 9.52217
R1984 VDPWR.n1155 VDPWR.t5 9.52217
R1985 VDPWR.n1155 VDPWR.t239 9.52217
R1986 VDPWR.n1154 VDPWR.t13 9.52217
R1987 VDPWR.n1154 VDPWR.t7 9.52217
R1988 VDPWR.n1301 VDPWR.t56 9.52217
R1989 VDPWR.n1301 VDPWR.t505 9.52217
R1990 VDPWR.n1151 VDPWR.t127 9.52217
R1991 VDPWR.n1151 VDPWR.t54 9.52217
R1992 VDPWR.n1150 VDPWR.t232 9.52217
R1993 VDPWR.n1150 VDPWR.t492 9.52217
R1994 VDPWR.n1149 VDPWR.t490 9.52217
R1995 VDPWR.n1149 VDPWR.t383 9.52217
R1996 VDPWR.n1317 VDPWR.t299 9.52217
R1997 VDPWR.n1317 VDPWR.t263 9.52217
R1998 VDPWR.n1146 VDPWR.t595 9.52217
R1999 VDPWR.n1146 VDPWR.t50 9.52217
R2000 VDPWR.n1145 VDPWR.t161 9.52217
R2001 VDPWR.n1145 VDPWR.t602 9.52217
R2002 VDPWR.n1144 VDPWR.t224 9.52217
R2003 VDPWR.n1144 VDPWR.t133 9.52217
R2004 VDPWR.n998 VDPWR.t106 9.52217
R2005 VDPWR.n998 VDPWR.t213 9.52217
R2006 VDPWR.n995 VDPWR.t102 9.52217
R2007 VDPWR.n995 VDPWR.t582 9.52217
R2008 VDPWR.n1015 VDPWR.t235 9.52217
R2009 VDPWR.n1015 VDPWR.t97 9.52217
R2010 VDPWR.n991 VDPWR.t620 9.52217
R2011 VDPWR.n991 VDPWR.t38 9.52217
R2012 VDPWR.n1033 VDPWR.t192 9.52217
R2013 VDPWR.n1033 VDPWR.t230 9.52217
R2014 VDPWR.n987 VDPWR.t347 9.52217
R2015 VDPWR.n987 VDPWR.t228 9.52217
R2016 VDPWR.n1051 VDPWR.t585 9.52217
R2017 VDPWR.n1051 VDPWR.t563 9.52217
R2018 VDPWR.n983 VDPWR.t63 9.52217
R2019 VDPWR.n983 VDPWR.t565 9.52217
R2020 VDPWR.n1069 VDPWR.t155 9.52217
R2021 VDPWR.n1069 VDPWR.t201 9.52217
R2022 VDPWR.n979 VDPWR.t539 9.52217
R2023 VDPWR.n979 VDPWR.t69 9.52217
R2024 VDPWR.n1087 VDPWR.t402 9.52217
R2025 VDPWR.n1087 VDPWR.t336 9.52217
R2026 VDPWR.n975 VDPWR.t537 9.52217
R2027 VDPWR.n975 VDPWR.t338 9.52217
R2028 VDPWR.n1105 VDPWR.t511 9.52217
R2029 VDPWR.n1105 VDPWR.t345 9.52217
R2030 VDPWR.n971 VDPWR.t513 9.52217
R2031 VDPWR.n971 VDPWR.t573 9.52217
R2032 VDPWR.n1123 VDPWR.t41 9.52217
R2033 VDPWR.n1123 VDPWR.t117 9.52217
R2034 VDPWR.n967 VDPWR.t318 9.52217
R2035 VDPWR.n967 VDPWR.t395 9.52217
R2036 VDPWR.n1391 VDPWR.t159 9.52217
R2037 VDPWR.n1391 VDPWR.t526 9.52217
R2038 VDPWR.n205 VDPWR.t222 9.52217
R2039 VDPWR.n205 VDPWR.t149 9.52217
R2040 VDPWR.n194 VDPWR.t593 9.52217
R2041 VDPWR.n194 VDPWR.t342 9.52217
R2042 VDPWR.n229 VDPWR.t266 9.52217
R2043 VDPWR.n229 VDPWR.t358 9.52217
R2044 VDPWR.n218 VDPWR.t95 9.52217
R2045 VDPWR.n218 VDPWR.t406 9.52217
R2046 VDPWR.n253 VDPWR.t79 9.52217
R2047 VDPWR.n253 VDPWR.t52 9.52217
R2048 VDPWR.n242 VDPWR.t259 9.52217
R2049 VDPWR.n242 VDPWR.t257 9.52217
R2050 VDPWR.n277 VDPWR.t555 9.52217
R2051 VDPWR.n277 VDPWR.t275 9.52217
R2052 VDPWR.n266 VDPWR.t245 9.52217
R2053 VDPWR.n266 VDPWR.t356 9.52217
R2054 VDPWR.n301 VDPWR.t124 9.52217
R2055 VDPWR.n301 VDPWR.t515 9.52217
R2056 VDPWR.n290 VDPWR.t203 9.52217
R2057 VDPWR.n290 VDPWR.t413 9.52217
R2058 VDPWR.n325 VDPWR.t421 9.52217
R2059 VDPWR.n325 VDPWR.t436 9.52217
R2060 VDPWR.n314 VDPWR.t509 9.52217
R2061 VDPWR.n314 VDPWR.t352 9.52217
R2062 VDPWR.n34 VDPWR.t450 9.52217
R2063 VDPWR.n34 VDPWR.t424 9.52217
R2064 VDPWR.n23 VDPWR.t547 9.52217
R2065 VDPWR.n23 VDPWR.t278 9.52217
R2066 VDPWR.n58 VDPWR.t418 9.52217
R2067 VDPWR.n58 VDPWR.t433 9.52217
R2068 VDPWR.n47 VDPWR.t612 9.52217
R2069 VDPWR.n47 VDPWR.t610 9.52217
R2070 VDPWR.n1540 VDPWR.t88 9.39094
R2071 VDPWR.n519 VDPWR.n518 8.66346
R2072 VDPWR.n156 VDPWR.n155 8.66346
R2073 VDPWR.n498 VDPWR.n497 7.70883
R2074 VDPWR.n509 VDPWR.n508 7.70883
R2075 VDPWR.n135 VDPWR.n134 7.70883
R2076 VDPWR.n146 VDPWR.n145 7.70883
R2077 VDPWR.n530 VDPWR.n529 7.4066
R2078 VDPWR.n1572 VDPWR.n1571 7.4066
R2079 VDPWR.n498 VDPWR.n179 6.57828
R2080 VDPWR.n509 VDPWR.n173 6.57828
R2081 VDPWR.n135 VDPWR.n8 6.57828
R2082 VDPWR.n146 VDPWR.n2 6.57828
R2083 VDPWR.n1009 VDPWR.n1007 5.44168
R2084 VDPWR.n1007 VDPWR.n1006 5.44168
R2085 VDPWR.n1027 VDPWR.n1025 5.44168
R2086 VDPWR.n1025 VDPWR.n1024 5.44168
R2087 VDPWR.n1045 VDPWR.n1043 5.44168
R2088 VDPWR.n1043 VDPWR.n1042 5.44168
R2089 VDPWR.n1063 VDPWR.n1061 5.44168
R2090 VDPWR.n1061 VDPWR.n1060 5.44168
R2091 VDPWR.n1081 VDPWR.n1079 5.44168
R2092 VDPWR.n1079 VDPWR.n1078 5.44168
R2093 VDPWR.n1099 VDPWR.n1097 5.44168
R2094 VDPWR.n1097 VDPWR.n1096 5.44168
R2095 VDPWR.n1117 VDPWR.n1115 5.44168
R2096 VDPWR.n1115 VDPWR.n1114 5.44168
R2097 VDPWR.n1135 VDPWR.n1133 5.44168
R2098 VDPWR.n1133 VDPWR.n1132 5.44168
R2099 VDPWR.n496 VDPWR.n495 5.33119
R2100 VDPWR.n133 VDPWR.n132 5.33119
R2101 VDPWR.n507 VDPWR.n506 5.31424
R2102 VDPWR.n144 VDPWR.n143 5.31424
R2103 VDPWR.n1199 VDPWR.n1189 5.0005
R2104 VDPWR.n1404 VDPWR.n1389 5.0005
R2105 VDPWR.n1566 VDPWR.n1334 4.63898
R2106 VDPWR.n580 VDPWR.n579 4.40526
R2107 VDPWR.n597 VDPWR.n596 4.40526
R2108 VDPWR.n614 VDPWR.n613 4.40526
R2109 VDPWR.n631 VDPWR.n630 4.40526
R2110 VDPWR.n648 VDPWR.n647 4.40526
R2111 VDPWR.n665 VDPWR.n664 4.40526
R2112 VDPWR.n682 VDPWR.n681 4.40526
R2113 VDPWR.n699 VDPWR.n698 4.40526
R2114 VDPWR.n1566 VDPWR.n1565 4.29701
R2115 VDPWR.n1198 VDPWR.n1196 3.72599
R2116 VDPWR.n1214 VDPWR.n1213 3.72599
R2117 VDPWR.n1230 VDPWR.n1229 3.72599
R2118 VDPWR.n1246 VDPWR.n1245 3.72599
R2119 VDPWR.n1262 VDPWR.n1261 3.72599
R2120 VDPWR.n1278 VDPWR.n1277 3.72599
R2121 VDPWR.n1294 VDPWR.n1293 3.72599
R2122 VDPWR.n1310 VDPWR.n1309 3.72599
R2123 VDPWR.n1326 VDPWR.n1325 3.72599
R2124 VDPWR.n1403 VDPWR.n1397 3.72599
R2125 VDPWR.n1399 VDPWR.n1398 3.72599
R2126 VDPWR.n1431 VDPWR.n1430 3.72599
R2127 VDPWR.n1425 VDPWR.n1424 3.72599
R2128 VDPWR.n1459 VDPWR.n1458 3.72599
R2129 VDPWR.n1453 VDPWR.n1452 3.72599
R2130 VDPWR.n1483 VDPWR.n1482 3.72599
R2131 VDPWR.n1568 VDPWR.n1567 3.19848
R2132 VDPWR.n1568 VDPWR.n535 3.17204
R2133 VDPWR.n357 VDPWR.n356 3.13979
R2134 VDPWR.n124 VDPWR.n123 3.13979
R2135 VDPWR.n90 VDPWR.n89 3.13979
R2136 VDPWR.n1141 VDPWR 2.86795
R2137 VDPWR.n863 VDPWR.t18 2.77153
R2138 VDPWR.n1000 VDPWR.n999 2.53478
R2139 VDPWR.n1007 VDPWR.n1002 2.35344
R2140 VDPWR.n1025 VDPWR.n1020 2.35344
R2141 VDPWR.n1043 VDPWR.n1038 2.35344
R2142 VDPWR.n1061 VDPWR.n1056 2.35344
R2143 VDPWR.n1079 VDPWR.n1074 2.35344
R2144 VDPWR.n1097 VDPWR.n1092 2.35344
R2145 VDPWR.n1115 VDPWR.n1110 2.35344
R2146 VDPWR.n1133 VDPWR.n1128 2.35344
R2147 VDPWR.n1536 VDPWR.n1535 2.3255
R2148 VDPWR.n1530 VDPWR.n1511 2.3255
R2149 VDPWR.n870 VDPWR.n869 2.3255
R2150 VDPWR.n873 VDPWR.n872 2.3255
R2151 VDPWR.n877 VDPWR.n876 2.3255
R2152 VDPWR.n880 VDPWR.n879 2.3255
R2153 VDPWR.n884 VDPWR.n883 2.3255
R2154 VDPWR.n887 VDPWR.n886 2.3255
R2155 VDPWR.n891 VDPWR.n890 2.3255
R2156 VDPWR.n894 VDPWR.n893 2.3255
R2157 VDPWR.n898 VDPWR.n897 2.3255
R2158 VDPWR.n901 VDPWR.n900 2.3255
R2159 VDPWR.n905 VDPWR.n904 2.3255
R2160 VDPWR.n908 VDPWR.n907 2.3255
R2161 VDPWR.n912 VDPWR.n911 2.3255
R2162 VDPWR.n915 VDPWR.n914 2.3255
R2163 VDPWR.n919 VDPWR.n918 2.3255
R2164 VDPWR.n922 VDPWR.n921 2.3255
R2165 VDPWR.n926 VDPWR.n925 2.3255
R2166 VDPWR.n929 VDPWR.n928 2.3255
R2167 VDPWR.n933 VDPWR.n932 2.3255
R2168 VDPWR.n936 VDPWR.n935 2.3255
R2169 VDPWR.n940 VDPWR.n939 2.3255
R2170 VDPWR.n943 VDPWR.n942 2.3255
R2171 VDPWR.n947 VDPWR.n946 2.3255
R2172 VDPWR.n950 VDPWR.n949 2.3255
R2173 VDPWR.n954 VDPWR.n953 2.3255
R2174 VDPWR.n957 VDPWR.n956 2.3255
R2175 VDPWR.n961 VDPWR.n960 2.3255
R2176 VDPWR.n964 VDPWR.n963 2.3255
R2177 VDPWR.n1546 VDPWR.n1545 2.3255
R2178 VDPWR.n1549 VDPWR.n1548 2.3255
R2179 VDPWR.n1553 VDPWR.n1552 2.3255
R2180 VDPWR.n1556 VDPWR.n1555 2.3255
R2181 VDPWR.n1560 VDPWR.n1559 2.3255
R2182 VDPWR.n1563 VDPWR.n1562 2.3255
R2183 VDPWR.n522 VDPWR.n521 2.3255
R2184 VDPWR.n349 VDPWR.n348 2.3255
R2185 VDPWR.n344 VDPWR.n343 2.3255
R2186 VDPWR.n383 VDPWR.n382 2.3255
R2187 VDPWR.n378 VDPWR.n377 2.3255
R2188 VDPWR.n409 VDPWR.n408 2.3255
R2189 VDPWR.n404 VDPWR.n403 2.3255
R2190 VDPWR.n435 VDPWR.n434 2.3255
R2191 VDPWR.n430 VDPWR.n429 2.3255
R2192 VDPWR.n461 VDPWR.n460 2.3255
R2193 VDPWR.n456 VDPWR.n455 2.3255
R2194 VDPWR.n487 VDPWR.n486 2.3255
R2195 VDPWR.n482 VDPWR.n481 2.3255
R2196 VDPWR.n159 VDPWR.n158 2.3255
R2197 VDPWR.n82 VDPWR.n81 2.3255
R2198 VDPWR.n77 VDPWR.n76 2.3255
R2199 VDPWR.n116 VDPWR.n115 2.3255
R2200 VDPWR.n111 VDPWR.n110 2.3255
R2201 VDPWR.n1011 VDPWR.n996 2.29581
R2202 VDPWR.n1014 VDPWR.n994 2.29581
R2203 VDPWR.n1018 VDPWR.n1017 2.29581
R2204 VDPWR.n1029 VDPWR.n992 2.29581
R2205 VDPWR.n1032 VDPWR.n990 2.29581
R2206 VDPWR.n1036 VDPWR.n1035 2.29581
R2207 VDPWR.n1047 VDPWR.n988 2.29581
R2208 VDPWR.n1050 VDPWR.n986 2.29581
R2209 VDPWR.n1054 VDPWR.n1053 2.29581
R2210 VDPWR.n1065 VDPWR.n984 2.29581
R2211 VDPWR.n1068 VDPWR.n982 2.29581
R2212 VDPWR.n1072 VDPWR.n1071 2.29581
R2213 VDPWR.n1083 VDPWR.n980 2.29581
R2214 VDPWR.n1086 VDPWR.n978 2.29581
R2215 VDPWR.n1090 VDPWR.n1089 2.29581
R2216 VDPWR.n1101 VDPWR.n976 2.29581
R2217 VDPWR.n1104 VDPWR.n974 2.29581
R2218 VDPWR.n1108 VDPWR.n1107 2.29581
R2219 VDPWR.n1119 VDPWR.n972 2.29581
R2220 VDPWR.n1122 VDPWR.n970 2.29581
R2221 VDPWR.n1126 VDPWR.n1125 2.29581
R2222 VDPWR.n1137 VDPWR.n968 2.29581
R2223 VDPWR.n1140 VDPWR.n966 2.29581
R2224 VDPWR.n359 VDPWR.n358 2.2505
R2225 VDPWR.n92 VDPWR.n91 2.2505
R2226 VDPWR.n126 VDPWR.n125 2.2505
R2227 VDPWR.n523 VDPWR.n514 2.2281
R2228 VDPWR.n160 VDPWR.n151 2.2281
R2229 VDPWR.n1193 VDPWR.n1192 2.1858
R2230 VDPWR.n520 VDPWR.n515 2.17472
R2231 VDPWR.n157 VDPWR.n152 2.17472
R2232 VDPWR.n1575 VDPWR.n1574 2.17342
R2233 VDPWR.n1570 VDPWR.n1569 2.17342
R2234 VDPWR.n1533 VDPWR.n1532 2.16821
R2235 VDPWR.n1538 VDPWR.n1528 2.16821
R2236 VDPWR.n1543 VDPWR.n1542 2.16821
R2237 VDPWR.n73 VDPWR.n44 2.16821
R2238 VDPWR.n591 VDPWR.n590 2.122
R2239 VDPWR.n608 VDPWR.n607 2.122
R2240 VDPWR.n625 VDPWR.n624 2.122
R2241 VDPWR.n642 VDPWR.n641 2.122
R2242 VDPWR.n659 VDPWR.n658 2.122
R2243 VDPWR.n676 VDPWR.n675 2.122
R2244 VDPWR.n693 VDPWR.n692 2.122
R2245 VDPWR.n710 VDPWR.n709 2.122
R2246 VDPWR.t16 VDPWR.t76 2.08383
R2247 VDPWR.t0 VDPWR.t165 2.08383
R2248 VDPWR.t461 VDPWR.t2 2.07474
R2249 VDPWR.t474 VDPWR.t414 2.07474
R2250 VDPWR.n1394 VDPWR.n1393 2.0647
R2251 VDPWR.n1564 VDPWR.n1490 2.04321
R2252 VDPWR.n1496 VDPWR.n1493 2.04321
R2253 VDPWR.n1557 VDPWR.n1497 2.04321
R2254 VDPWR.n1503 VDPWR.n1500 2.04321
R2255 VDPWR.n1550 VDPWR.n1504 2.04321
R2256 VDPWR.n1510 VDPWR.n1507 2.04321
R2257 VDPWR.n866 VDPWR.n805 2.04321
R2258 VDPWR.n965 VDPWR.n711 2.04321
R2259 VDPWR.n717 VDPWR.n714 2.04321
R2260 VDPWR.n958 VDPWR.n718 2.04321
R2261 VDPWR.n724 VDPWR.n721 2.04321
R2262 VDPWR.n951 VDPWR.n725 2.04321
R2263 VDPWR.n731 VDPWR.n728 2.04321
R2264 VDPWR.n944 VDPWR.n732 2.04321
R2265 VDPWR.n738 VDPWR.n735 2.04321
R2266 VDPWR.n937 VDPWR.n739 2.04321
R2267 VDPWR.n745 VDPWR.n742 2.04321
R2268 VDPWR.n930 VDPWR.n746 2.04321
R2269 VDPWR.n752 VDPWR.n749 2.04321
R2270 VDPWR.n923 VDPWR.n753 2.04321
R2271 VDPWR.n759 VDPWR.n756 2.04321
R2272 VDPWR.n916 VDPWR.n760 2.04321
R2273 VDPWR.n766 VDPWR.n763 2.04321
R2274 VDPWR.n909 VDPWR.n767 2.04321
R2275 VDPWR.n773 VDPWR.n770 2.04321
R2276 VDPWR.n902 VDPWR.n774 2.04321
R2277 VDPWR.n780 VDPWR.n777 2.04321
R2278 VDPWR.n895 VDPWR.n781 2.04321
R2279 VDPWR.n787 VDPWR.n784 2.04321
R2280 VDPWR.n888 VDPWR.n788 2.04321
R2281 VDPWR.n794 VDPWR.n791 2.04321
R2282 VDPWR.n881 VDPWR.n795 2.04321
R2283 VDPWR.n801 VDPWR.n798 2.04321
R2284 VDPWR.n874 VDPWR.n802 2.04321
R2285 VDPWR.n867 VDPWR.n865 2.04321
R2286 VDPWR.n479 VDPWR.n192 2.04321
R2287 VDPWR.n478 VDPWR.n191 2.04321
R2288 VDPWR.n185 VDPWR.n184 2.04321
R2289 VDPWR.n489 VDPWR.n183 2.04321
R2290 VDPWR.n453 VDPWR.n216 2.04321
R2291 VDPWR.n452 VDPWR.n215 2.04321
R2292 VDPWR.n209 VDPWR.n208 2.04321
R2293 VDPWR.n463 VDPWR.n207 2.04321
R2294 VDPWR.n427 VDPWR.n240 2.04321
R2295 VDPWR.n426 VDPWR.n239 2.04321
R2296 VDPWR.n233 VDPWR.n232 2.04321
R2297 VDPWR.n437 VDPWR.n231 2.04321
R2298 VDPWR.n401 VDPWR.n264 2.04321
R2299 VDPWR.n400 VDPWR.n263 2.04321
R2300 VDPWR.n257 VDPWR.n256 2.04321
R2301 VDPWR.n411 VDPWR.n255 2.04321
R2302 VDPWR.n375 VDPWR.n288 2.04321
R2303 VDPWR.n374 VDPWR.n287 2.04321
R2304 VDPWR.n281 VDPWR.n280 2.04321
R2305 VDPWR.n385 VDPWR.n279 2.04321
R2306 VDPWR.n341 VDPWR.n312 2.04321
R2307 VDPWR.n340 VDPWR.n311 2.04321
R2308 VDPWR.n305 VDPWR.n304 2.04321
R2309 VDPWR.n351 VDPWR.n303 2.04321
R2310 VDPWR.n108 VDPWR.n21 2.04321
R2311 VDPWR.n107 VDPWR.n20 2.04321
R2312 VDPWR.n14 VDPWR.n13 2.04321
R2313 VDPWR.n118 VDPWR.n12 2.04321
R2314 VDPWR.n74 VDPWR.n45 2.04321
R2315 VDPWR.n84 VDPWR.n36 2.04321
R2316 VDPWR.n38 VDPWR.n37 2.04321
R2317 VDPWR.n527 VDPWR.n526 2.0406
R2318 VDPWR.n535 VDPWR.n167 2.0406
R2319 VDPWR.n525 VDPWR.n170 1.99827
R2320 VDPWR.n1006 VDPWR.n1005 1.97967
R2321 VDPWR.n1024 VDPWR.n1023 1.97967
R2322 VDPWR.n1042 VDPWR.n1041 1.97967
R2323 VDPWR.n1060 VDPWR.n1059 1.97967
R2324 VDPWR.n1078 VDPWR.n1077 1.97967
R2325 VDPWR.n1096 VDPWR.n1095 1.97967
R2326 VDPWR.n1114 VDPWR.n1113 1.97967
R2327 VDPWR.n1132 VDPWR.n1131 1.97967
R2328 VDPWR VDPWR.n324 1.97234
R2329 VDPWR VDPWR.n57 1.97234
R2330 VDPWR.n493 VDPWR.n492 1.96588
R2331 VDPWR.n501 VDPWR.n177 1.96588
R2332 VDPWR.n504 VDPWR.n503 1.96588
R2333 VDPWR.n512 VDPWR.n171 1.96588
R2334 VDPWR.n130 VDPWR.n129 1.96588
R2335 VDPWR.n138 VDPWR.n6 1.96588
R2336 VDPWR.n141 VDPWR.n140 1.96588
R2337 VDPWR.n149 VDPWR.n0 1.96588
R2338 VDPWR.n468 VDPWR.n201 1.96583
R2339 VDPWR.n464 VDPWR.n204 1.96583
R2340 VDPWR.n197 VDPWR.n196 1.96583
R2341 VDPWR.n477 VDPWR.n193 1.96583
R2342 VDPWR.n442 VDPWR.n225 1.96583
R2343 VDPWR.n438 VDPWR.n228 1.96583
R2344 VDPWR.n221 VDPWR.n220 1.96583
R2345 VDPWR.n451 VDPWR.n217 1.96583
R2346 VDPWR.n416 VDPWR.n249 1.96583
R2347 VDPWR.n412 VDPWR.n252 1.96583
R2348 VDPWR.n245 VDPWR.n244 1.96583
R2349 VDPWR.n425 VDPWR.n241 1.96583
R2350 VDPWR.n390 VDPWR.n273 1.96583
R2351 VDPWR.n386 VDPWR.n276 1.96583
R2352 VDPWR.n269 VDPWR.n268 1.96583
R2353 VDPWR.n399 VDPWR.n265 1.96583
R2354 VDPWR.n364 VDPWR.n297 1.96583
R2355 VDPWR.n360 VDPWR.n300 1.96583
R2356 VDPWR.n293 VDPWR.n292 1.96583
R2357 VDPWR.n373 VDPWR.n289 1.96583
R2358 VDPWR.n330 VDPWR.n321 1.96583
R2359 VDPWR.n317 VDPWR.n316 1.96583
R2360 VDPWR.n339 VDPWR.n313 1.96583
R2361 VDPWR.n97 VDPWR.n30 1.96583
R2362 VDPWR.n93 VDPWR.n33 1.96583
R2363 VDPWR.n26 VDPWR.n25 1.96583
R2364 VDPWR.n106 VDPWR.n22 1.96583
R2365 VDPWR.n63 VDPWR.n54 1.96583
R2366 VDPWR.n50 VDPWR.n49 1.96583
R2367 VDPWR.n72 VDPWR.n46 1.96583
R2368 VDPWR.n1204 VDPWR.n1183 1.9397
R2369 VDPWR.n1208 VDPWR.n1207 1.9397
R2370 VDPWR.n1220 VDPWR.n1178 1.9397
R2371 VDPWR.n1224 VDPWR.n1223 1.9397
R2372 VDPWR.n1236 VDPWR.n1173 1.9397
R2373 VDPWR.n1240 VDPWR.n1239 1.9397
R2374 VDPWR.n1252 VDPWR.n1168 1.9397
R2375 VDPWR.n1256 VDPWR.n1255 1.9397
R2376 VDPWR.n1268 VDPWR.n1163 1.9397
R2377 VDPWR.n1272 VDPWR.n1271 1.9397
R2378 VDPWR.n1284 VDPWR.n1158 1.9397
R2379 VDPWR.n1288 VDPWR.n1287 1.9397
R2380 VDPWR.n1300 VDPWR.n1153 1.9397
R2381 VDPWR.n1304 VDPWR.n1303 1.9397
R2382 VDPWR.n1316 VDPWR.n1148 1.9397
R2383 VDPWR.n1320 VDPWR.n1319 1.9397
R2384 VDPWR.n1332 VDPWR.n1143 1.9397
R2385 VDPWR.n1409 VDPWR.n1383 1.9397
R2386 VDPWR.n1410 VDPWR.n1379 1.9397
R2387 VDPWR.n1419 VDPWR.n1378 1.9397
R2388 VDPWR.n1377 VDPWR.n1372 1.9397
R2389 VDPWR.n1437 VDPWR.n1367 1.9397
R2390 VDPWR.n1438 VDPWR.n1363 1.9397
R2391 VDPWR.n1447 VDPWR.n1362 1.9397
R2392 VDPWR.n1361 VDPWR.n1356 1.9397
R2393 VDPWR.n1465 VDPWR.n1351 1.9397
R2394 VDPWR.n1466 VDPWR.n1347 1.9397
R2395 VDPWR.n1475 VDPWR.n1346 1.9397
R2396 VDPWR.n1345 VDPWR.n1340 1.9397
R2397 VDPWR.n1489 VDPWR.n1335 1.9397
R2398 VDPWR.n533 VDPWR.n532 1.8605
R2399 VDPWR.n165 VDPWR.n163 1.8605
R2400 VDPWR.n181 VDPWR.n178 1.54255
R2401 VDPWR.n175 VDPWR.n172 1.54255
R2402 VDPWR.n10 VDPWR.n7 1.54255
R2403 VDPWR.n4 VDPWR.n1 1.54255
R2404 VDPWR.n1207 VDPWR.n1204 1.52654
R2405 VDPWR.n1223 VDPWR.n1220 1.52654
R2406 VDPWR.n1239 VDPWR.n1236 1.52654
R2407 VDPWR.n1255 VDPWR.n1252 1.52654
R2408 VDPWR.n1271 VDPWR.n1268 1.52654
R2409 VDPWR.n1287 VDPWR.n1284 1.52654
R2410 VDPWR.n1303 VDPWR.n1300 1.52654
R2411 VDPWR.n1319 VDPWR.n1316 1.52654
R2412 VDPWR.n705 VDPWR.n701 1.51949
R2413 VDPWR.n688 VDPWR.n684 1.51949
R2414 VDPWR.n671 VDPWR.n667 1.51949
R2415 VDPWR.n654 VDPWR.n650 1.51949
R2416 VDPWR.n637 VDPWR.n633 1.51949
R2417 VDPWR.n620 VDPWR.n616 1.51949
R2418 VDPWR.n603 VDPWR.n599 1.51949
R2419 VDPWR.n586 VDPWR.n582 1.51949
R2420 VDPWR.n1569 VDPWR.n1568 1.45922
R2421 VDPWR.n1333 VDPWR.n1142 1.39972
R2422 VDPWR.n129 VDPWR 1.37724
R2423 VDPWR.n337 VDPWR.n336 1.32907
R2424 VDPWR.n329 VDPWR.n328 1.32907
R2425 VDPWR.n371 VDPWR.n370 1.32907
R2426 VDPWR.n363 VDPWR.n362 1.32907
R2427 VDPWR.n397 VDPWR.n396 1.32907
R2428 VDPWR.n389 VDPWR.n388 1.32907
R2429 VDPWR.n423 VDPWR.n422 1.32907
R2430 VDPWR.n415 VDPWR.n414 1.32907
R2431 VDPWR.n449 VDPWR.n448 1.32907
R2432 VDPWR.n441 VDPWR.n440 1.32907
R2433 VDPWR.n475 VDPWR.n474 1.32907
R2434 VDPWR.n467 VDPWR.n466 1.32907
R2435 VDPWR.n70 VDPWR.n69 1.32907
R2436 VDPWR.n62 VDPWR.n61 1.32907
R2437 VDPWR.n104 VDPWR.n103 1.32907
R2438 VDPWR.n96 VDPWR.n95 1.32907
R2439 VDPWR.n356 VDPWR 1.24128
R2440 VDPWR.n123 VDPWR 1.24128
R2441 VDPWR.n89 VDPWR 1.24128
R2442 VDPWR.n492 VDPWR 1.23314
R2443 VDPWR.n465 VDPWR.n206 1.21789
R2444 VDPWR.n476 VDPWR.n195 1.21789
R2445 VDPWR.n439 VDPWR.n230 1.21789
R2446 VDPWR.n450 VDPWR.n219 1.21789
R2447 VDPWR.n413 VDPWR.n254 1.21789
R2448 VDPWR.n424 VDPWR.n243 1.21789
R2449 VDPWR.n387 VDPWR.n278 1.21789
R2450 VDPWR.n398 VDPWR.n267 1.21789
R2451 VDPWR.n361 VDPWR.n302 1.21789
R2452 VDPWR.n372 VDPWR.n291 1.21789
R2453 VDPWR.n327 VDPWR.n326 1.21789
R2454 VDPWR.n338 VDPWR.n315 1.21789
R2455 VDPWR.n94 VDPWR.n35 1.21789
R2456 VDPWR.n105 VDPWR.n24 1.21789
R2457 VDPWR.n60 VDPWR.n59 1.21789
R2458 VDPWR.n71 VDPWR.n48 1.21789
R2459 VDPWR.n1216 VDPWR.n1215 1.21332
R2460 VDPWR.n1232 VDPWR.n1231 1.21332
R2461 VDPWR.n1248 VDPWR.n1247 1.21332
R2462 VDPWR.n1264 VDPWR.n1263 1.21332
R2463 VDPWR.n1280 VDPWR.n1279 1.21332
R2464 VDPWR.n1296 VDPWR.n1295 1.21332
R2465 VDPWR.n1312 VDPWR.n1311 1.21332
R2466 VDPWR.n1328 VDPWR.n1327 1.21332
R2467 VDPWR.n1418 VDPWR.n1380 1.21332
R2468 VDPWR.n1433 VDPWR.n1432 1.21332
R2469 VDPWR.n1446 VDPWR.n1364 1.21332
R2470 VDPWR.n1461 VDPWR.n1460 1.21332
R2471 VDPWR.n1474 VDPWR.n1348 1.21332
R2472 VDPWR.n1485 VDPWR.n1484 1.21332
R2473 VDPWR.n354 VDPWR.n353 1.09595
R2474 VDPWR.n121 VDPWR.n120 1.09595
R2475 VDPWR.n87 VDPWR.n86 1.09595
R2476 VDPWR.n592 VDPWR 1.04243
R2477 VDPWR.n609 VDPWR 1.04243
R2478 VDPWR.n626 VDPWR 1.04243
R2479 VDPWR.n643 VDPWR 1.04243
R2480 VDPWR.n660 VDPWR 1.04243
R2481 VDPWR.n677 VDPWR 1.04243
R2482 VDPWR.n694 VDPWR 1.04243
R2483 VDPWR.n1141 VDPWR.n965 0.948417
R2484 VDPWR.n572 VDPWR.n571 0.832022
R2485 VDPWR.n567 VDPWR.n566 0.832022
R2486 VDPWR.n562 VDPWR.n561 0.832022
R2487 VDPWR.n557 VDPWR.n556 0.832022
R2488 VDPWR.n552 VDPWR.n551 0.832022
R2489 VDPWR.n547 VDPWR.n546 0.832022
R2490 VDPWR.n542 VDPWR.n541 0.832022
R2491 VDPWR.n537 VDPWR.n536 0.832022
R2492 VDPWR VDPWR.n1332 0.813
R2493 VDPWR.n358 VDPWR.n357 0.8005
R2494 VDPWR.n91 VDPWR.n90 0.795143
R2495 VDPWR.n125 VDPWR.n124 0.777286
R2496 VDPWR.n127 VDPWR 0.7505
R2497 VDPWR.n1567 VDPWR.n1566 0.68153
R2498 VDPWR.n1017 VDPWR 0.669618
R2499 VDPWR.n1035 VDPWR 0.669618
R2500 VDPWR.n1053 VDPWR 0.669618
R2501 VDPWR.n1071 VDPWR 0.669618
R2502 VDPWR.n1089 VDPWR 0.669618
R2503 VDPWR.n1107 VDPWR 0.669618
R2504 VDPWR.n1125 VDPWR 0.669618
R2505 VDPWR.n524 VDPWR.n513 0.6555
R2506 VDPWR.n161 VDPWR.n150 0.6555
R2507 VDPWR.n576 VDPWR.n574 0.629553
R2508 VDPWR.n1329 VDPWR.n1328 0.6205
R2509 VDPWR.n1313 VDPWR.n1312 0.6205
R2510 VDPWR.n1297 VDPWR.n1296 0.6205
R2511 VDPWR.n1281 VDPWR.n1280 0.6205
R2512 VDPWR.n1265 VDPWR.n1264 0.6205
R2513 VDPWR.n1249 VDPWR.n1248 0.6205
R2514 VDPWR.n1233 VDPWR.n1232 0.6205
R2515 VDPWR.n1217 VDPWR.n1216 0.6205
R2516 VDPWR.n1201 VDPWR.n1200 0.6205
R2517 VDPWR.n1486 VDPWR.n1485 0.6205
R2518 VDPWR.n1474 VDPWR.n1473 0.6205
R2519 VDPWR.n1462 VDPWR.n1461 0.6205
R2520 VDPWR.n1446 VDPWR.n1445 0.6205
R2521 VDPWR.n1434 VDPWR.n1433 0.6205
R2522 VDPWR.n1418 VDPWR.n1417 0.6205
R2523 VDPWR.n1406 VDPWR.n1405 0.6205
R2524 VDPWR.n574 VDPWR.n573 0.61463
R2525 VDPWR.n569 VDPWR.n568 0.61463
R2526 VDPWR.n564 VDPWR.n563 0.61463
R2527 VDPWR.n559 VDPWR.n558 0.61463
R2528 VDPWR.n554 VDPWR.n553 0.61463
R2529 VDPWR.n549 VDPWR.n548 0.61463
R2530 VDPWR.n544 VDPWR.n543 0.61463
R2531 VDPWR.n539 VDPWR.n538 0.61463
R2532 VDPWR.n1575 VDPWR.n161 0.60099
R2533 VDPWR.n1136 VDPWR.n1135 0.58175
R2534 VDPWR.n1118 VDPWR.n1117 0.58175
R2535 VDPWR.n1100 VDPWR.n1099 0.58175
R2536 VDPWR.n1082 VDPWR.n1081 0.58175
R2537 VDPWR.n1064 VDPWR.n1063 0.58175
R2538 VDPWR.n1046 VDPWR.n1045 0.58175
R2539 VDPWR.n1028 VDPWR.n1027 0.58175
R2540 VDPWR.n1010 VDPWR.n1009 0.58175
R2541 VDPWR VDPWR.n385 0.568208
R2542 VDPWR VDPWR.n411 0.568208
R2543 VDPWR VDPWR.n437 0.568208
R2544 VDPWR VDPWR.n463 0.568208
R2545 VDPWR.n1200 VDPWR.n1188 0.533833
R2546 VDPWR.n1405 VDPWR.n1388 0.533833
R2547 VDPWR.n525 VDPWR.n524 0.517657
R2548 VDPWR.n513 VDPWR 0.472722
R2549 VDPWR.n150 VDPWR 0.472722
R2550 VDPWR.n503 VDPWR 0.453625
R2551 VDPWR.n140 VDPWR 0.453625
R2552 VDPWR.n340 VDPWR 0.432792
R2553 VDPWR.n374 VDPWR 0.432792
R2554 VDPWR.n400 VDPWR 0.432792
R2555 VDPWR.n426 VDPWR 0.432792
R2556 VDPWR.n452 VDPWR 0.432792
R2557 VDPWR.n478 VDPWR 0.432792
R2558 VDPWR.n107 VDPWR 0.432792
R2559 VDPWR.n321 VDPWR.n316 0.430188
R2560 VDPWR.n297 VDPWR.n292 0.430188
R2561 VDPWR.n273 VDPWR.n268 0.430188
R2562 VDPWR.n249 VDPWR.n244 0.430188
R2563 VDPWR.n225 VDPWR.n220 0.430188
R2564 VDPWR.n201 VDPWR.n196 0.430188
R2565 VDPWR.n54 VDPWR.n49 0.430188
R2566 VDPWR.n30 VDPWR.n25 0.430188
R2567 VDPWR.n510 VDPWR.n509 0.423227
R2568 VDPWR.n499 VDPWR.n498 0.423227
R2569 VDPWR.n147 VDPWR.n146 0.423227
R2570 VDPWR.n136 VDPWR.n135 0.423227
R2571 VDPWR.n356 VDPWR 0.402286
R2572 VDPWR.n123 VDPWR 0.402286
R2573 VDPWR.n89 VDPWR 0.402286
R2574 VDPWR.n73 VDPWR 0.401542
R2575 VDPWR.n1567 VDPWR 0.392832
R2576 VDPWR VDPWR.n359 0.389823
R2577 VDPWR VDPWR.n92 0.385917
R2578 VDPWR VDPWR.n591 0.3755
R2579 VDPWR VDPWR.n608 0.3755
R2580 VDPWR VDPWR.n625 0.3755
R2581 VDPWR VDPWR.n642 0.3755
R2582 VDPWR VDPWR.n659 0.3755
R2583 VDPWR VDPWR.n676 0.3755
R2584 VDPWR VDPWR.n693 0.3755
R2585 VDPWR VDPWR.n710 0.3755
R2586 VDPWR.n328 VDPWR.n321 0.359875
R2587 VDPWR.n337 VDPWR.n316 0.359875
R2588 VDPWR.n362 VDPWR.n297 0.359875
R2589 VDPWR.n371 VDPWR.n292 0.359875
R2590 VDPWR.n388 VDPWR.n273 0.359875
R2591 VDPWR.n397 VDPWR.n268 0.359875
R2592 VDPWR.n414 VDPWR.n249 0.359875
R2593 VDPWR.n423 VDPWR.n244 0.359875
R2594 VDPWR.n440 VDPWR.n225 0.359875
R2595 VDPWR.n449 VDPWR.n220 0.359875
R2596 VDPWR.n466 VDPWR.n201 0.359875
R2597 VDPWR.n475 VDPWR.n196 0.359875
R2598 VDPWR.n61 VDPWR.n54 0.359875
R2599 VDPWR.n70 VDPWR.n49 0.359875
R2600 VDPWR.n95 VDPWR.n30 0.359875
R2601 VDPWR.n104 VDPWR.n25 0.359875
R2602 VDPWR.n593 VDPWR.n592 0.358192
R2603 VDPWR.n610 VDPWR.n609 0.358192
R2604 VDPWR.n627 VDPWR.n626 0.358192
R2605 VDPWR.n644 VDPWR.n643 0.358192
R2606 VDPWR.n661 VDPWR.n660 0.358192
R2607 VDPWR.n678 VDPWR.n677 0.358192
R2608 VDPWR.n695 VDPWR.n694 0.358192
R2609 VDPWR.n490 VDPWR.n489 0.357271
R2610 VDPWR.n573 VDPWR.n572 0.353761
R2611 VDPWR.n568 VDPWR.n567 0.353761
R2612 VDPWR.n563 VDPWR.n562 0.353761
R2613 VDPWR.n558 VDPWR.n557 0.353761
R2614 VDPWR.n553 VDPWR.n552 0.353761
R2615 VDPWR.n548 VDPWR.n547 0.353761
R2616 VDPWR.n543 VDPWR.n542 0.353761
R2617 VDPWR.n538 VDPWR.n537 0.353761
R2618 VDPWR.n1142 VDPWR 0.350184
R2619 VDPWR.n490 VDPWR 0.333833
R2620 VDPWR.n999 VDPWR.n997 0.324029
R2621 VDPWR.n1013 VDPWR.n1012 0.324029
R2622 VDPWR.n1016 VDPWR.n993 0.324029
R2623 VDPWR.n1031 VDPWR.n1030 0.324029
R2624 VDPWR.n1034 VDPWR.n989 0.324029
R2625 VDPWR.n1049 VDPWR.n1048 0.324029
R2626 VDPWR.n1052 VDPWR.n985 0.324029
R2627 VDPWR.n1067 VDPWR.n1066 0.324029
R2628 VDPWR.n1070 VDPWR.n981 0.324029
R2629 VDPWR.n1085 VDPWR.n1084 0.324029
R2630 VDPWR.n1088 VDPWR.n977 0.324029
R2631 VDPWR.n1103 VDPWR.n1102 0.324029
R2632 VDPWR.n1106 VDPWR.n973 0.324029
R2633 VDPWR.n1121 VDPWR.n1120 0.324029
R2634 VDPWR.n1124 VDPWR.n969 0.324029
R2635 VDPWR.n1139 VDPWR.n1138 0.324029
R2636 VDPWR.n1142 VDPWR.n1141 0.274719
R2637 VDPWR.n592 VDPWR.n569 0.271861
R2638 VDPWR.n609 VDPWR.n564 0.271861
R2639 VDPWR.n626 VDPWR.n559 0.271861
R2640 VDPWR.n643 VDPWR.n554 0.271861
R2641 VDPWR.n660 VDPWR.n549 0.271861
R2642 VDPWR.n677 VDPWR.n544 0.271861
R2643 VDPWR.n694 VDPWR.n539 0.271861
R2644 VDPWR.n1201 VDPWR.n1187 0.253104
R2645 VDPWR.n1217 VDPWR.n1182 0.253104
R2646 VDPWR.n1233 VDPWR.n1177 0.253104
R2647 VDPWR.n1249 VDPWR.n1172 0.253104
R2648 VDPWR.n1265 VDPWR.n1167 0.253104
R2649 VDPWR.n1281 VDPWR.n1162 0.253104
R2650 VDPWR.n1297 VDPWR.n1157 0.253104
R2651 VDPWR.n1313 VDPWR.n1152 0.253104
R2652 VDPWR.n1329 VDPWR.n1147 0.253104
R2653 VDPWR.n1406 VDPWR.n1387 0.253104
R2654 VDPWR.n1417 VDPWR.n1412 0.253104
R2655 VDPWR.n1434 VDPWR.n1371 0.253104
R2656 VDPWR.n1445 VDPWR.n1440 0.253104
R2657 VDPWR.n1462 VDPWR.n1355 0.253104
R2658 VDPWR.n1473 VDPWR.n1468 0.253104
R2659 VDPWR.n1486 VDPWR.n1339 0.253104
R2660 VDPWR.n1009 VDPWR.n1008 0.25148
R2661 VDPWR.n1027 VDPWR.n1026 0.25148
R2662 VDPWR.n1045 VDPWR.n1044 0.25148
R2663 VDPWR.n1063 VDPWR.n1062 0.25148
R2664 VDPWR.n1081 VDPWR.n1080 0.25148
R2665 VDPWR.n1099 VDPWR.n1098 0.25148
R2666 VDPWR.n1117 VDPWR.n1116 0.25148
R2667 VDPWR.n1135 VDPWR.n1134 0.25148
R2668 VDPWR.n1204 VDPWR.n1203 0.246594
R2669 VDPWR.n1207 VDPWR.n1206 0.246594
R2670 VDPWR.n1220 VDPWR.n1219 0.246594
R2671 VDPWR.n1223 VDPWR.n1222 0.246594
R2672 VDPWR.n1236 VDPWR.n1235 0.246594
R2673 VDPWR.n1239 VDPWR.n1238 0.246594
R2674 VDPWR.n1252 VDPWR.n1251 0.246594
R2675 VDPWR.n1255 VDPWR.n1254 0.246594
R2676 VDPWR.n1268 VDPWR.n1267 0.246594
R2677 VDPWR.n1271 VDPWR.n1270 0.246594
R2678 VDPWR.n1284 VDPWR.n1283 0.246594
R2679 VDPWR.n1287 VDPWR.n1286 0.246594
R2680 VDPWR.n1300 VDPWR.n1299 0.246594
R2681 VDPWR.n1303 VDPWR.n1302 0.246594
R2682 VDPWR.n1316 VDPWR.n1315 0.246594
R2683 VDPWR.n1319 VDPWR.n1318 0.246594
R2684 VDPWR.n1332 VDPWR.n1331 0.246594
R2685 VDPWR.n1409 VDPWR.n1408 0.246594
R2686 VDPWR.n1411 VDPWR.n1410 0.246594
R2687 VDPWR.n1415 VDPWR.n1378 0.246594
R2688 VDPWR.n1377 VDPWR.n1376 0.246594
R2689 VDPWR.n1437 VDPWR.n1436 0.246594
R2690 VDPWR.n1439 VDPWR.n1438 0.246594
R2691 VDPWR.n1443 VDPWR.n1362 0.246594
R2692 VDPWR.n1361 VDPWR.n1360 0.246594
R2693 VDPWR.n1465 VDPWR.n1464 0.246594
R2694 VDPWR.n1467 VDPWR.n1466 0.246594
R2695 VDPWR.n1471 VDPWR.n1346 0.246594
R2696 VDPWR.n1345 VDPWR.n1344 0.246594
R2697 VDPWR.n1489 VDPWR.n1488 0.246594
R2698 VDPWR.n1202 VDPWR.n1201 0.242688
R2699 VDPWR.n1218 VDPWR.n1217 0.242688
R2700 VDPWR.n1234 VDPWR.n1233 0.242688
R2701 VDPWR.n1250 VDPWR.n1249 0.242688
R2702 VDPWR.n1266 VDPWR.n1265 0.242688
R2703 VDPWR.n1282 VDPWR.n1281 0.242688
R2704 VDPWR.n1298 VDPWR.n1297 0.242688
R2705 VDPWR.n1314 VDPWR.n1313 0.242688
R2706 VDPWR.n1330 VDPWR.n1329 0.242688
R2707 VDPWR.n1407 VDPWR.n1406 0.242688
R2708 VDPWR.n1417 VDPWR.n1416 0.242688
R2709 VDPWR.n1435 VDPWR.n1434 0.242688
R2710 VDPWR.n1445 VDPWR.n1444 0.242688
R2711 VDPWR.n1463 VDPWR.n1462 0.242688
R2712 VDPWR.n1473 VDPWR.n1472 0.242688
R2713 VDPWR.n1487 VDPWR.n1486 0.242688
R2714 VDPWR.n1565 VDPWR 0.240083
R2715 VDPWR.n1017 VDPWR.n1016 0.239471
R2716 VDPWR.n1035 VDPWR.n1034 0.239471
R2717 VDPWR.n1053 VDPWR.n1052 0.239471
R2718 VDPWR.n1071 VDPWR.n1070 0.239471
R2719 VDPWR.n1089 VDPWR.n1088 0.239471
R2720 VDPWR.n1107 VDPWR.n1106 0.239471
R2721 VDPWR.n1125 VDPWR.n1124 0.239471
R2722 VDPWR.n1014 VDPWR.n1013 0.232118
R2723 VDPWR.n1032 VDPWR.n1031 0.232118
R2724 VDPWR.n1050 VDPWR.n1049 0.232118
R2725 VDPWR.n1068 VDPWR.n1067 0.232118
R2726 VDPWR.n1086 VDPWR.n1085 0.232118
R2727 VDPWR.n1104 VDPWR.n1103 0.232118
R2728 VDPWR.n1122 VDPWR.n1121 0.232118
R2729 VDPWR.n1140 VDPWR.n1139 0.232118
R2730 VDPWR.n1192 VDPWR.n1187 0.229667
R2731 VDPWR.n1203 VDPWR.n1202 0.229667
R2732 VDPWR.n1206 VDPWR.n1182 0.229667
R2733 VDPWR.n1219 VDPWR.n1218 0.229667
R2734 VDPWR.n1222 VDPWR.n1177 0.229667
R2735 VDPWR.n1235 VDPWR.n1234 0.229667
R2736 VDPWR.n1238 VDPWR.n1172 0.229667
R2737 VDPWR.n1251 VDPWR.n1250 0.229667
R2738 VDPWR.n1254 VDPWR.n1167 0.229667
R2739 VDPWR.n1267 VDPWR.n1266 0.229667
R2740 VDPWR.n1270 VDPWR.n1162 0.229667
R2741 VDPWR.n1283 VDPWR.n1282 0.229667
R2742 VDPWR.n1286 VDPWR.n1157 0.229667
R2743 VDPWR.n1299 VDPWR.n1298 0.229667
R2744 VDPWR.n1302 VDPWR.n1152 0.229667
R2745 VDPWR.n1315 VDPWR.n1314 0.229667
R2746 VDPWR.n1318 VDPWR.n1147 0.229667
R2747 VDPWR.n1331 VDPWR.n1330 0.229667
R2748 VDPWR.n1408 VDPWR.n1407 0.229667
R2749 VDPWR.n1412 VDPWR.n1411 0.229667
R2750 VDPWR.n1416 VDPWR.n1415 0.229667
R2751 VDPWR.n1376 VDPWR.n1371 0.229667
R2752 VDPWR.n1436 VDPWR.n1435 0.229667
R2753 VDPWR.n1440 VDPWR.n1439 0.229667
R2754 VDPWR.n1444 VDPWR.n1443 0.229667
R2755 VDPWR.n1360 VDPWR.n1355 0.229667
R2756 VDPWR.n1464 VDPWR.n1463 0.229667
R2757 VDPWR.n1468 VDPWR.n1467 0.229667
R2758 VDPWR.n1472 VDPWR.n1471 0.229667
R2759 VDPWR.n1344 VDPWR.n1339 0.229667
R2760 VDPWR.n1488 VDPWR.n1487 0.229667
R2761 VDPWR.n328 VDPWR.n327 0.229667
R2762 VDPWR.n338 VDPWR.n337 0.229667
R2763 VDPWR.n362 VDPWR.n361 0.229667
R2764 VDPWR.n372 VDPWR.n371 0.229667
R2765 VDPWR.n388 VDPWR.n387 0.229667
R2766 VDPWR.n398 VDPWR.n397 0.229667
R2767 VDPWR.n414 VDPWR.n413 0.229667
R2768 VDPWR.n424 VDPWR.n423 0.229667
R2769 VDPWR.n440 VDPWR.n439 0.229667
R2770 VDPWR.n450 VDPWR.n449 0.229667
R2771 VDPWR.n466 VDPWR.n465 0.229667
R2772 VDPWR.n476 VDPWR.n475 0.229667
R2773 VDPWR.n61 VDPWR.n60 0.229667
R2774 VDPWR.n71 VDPWR.n70 0.229667
R2775 VDPWR.n95 VDPWR.n94 0.229667
R2776 VDPWR.n105 VDPWR.n104 0.229667
R2777 VDPWR.n524 VDPWR.n523 0.223
R2778 VDPWR.n161 VDPWR.n160 0.223
R2779 VDPWR.n1410 VDPWR.n1409 0.221854
R2780 VDPWR.n1378 VDPWR.n1377 0.221854
R2781 VDPWR.n1438 VDPWR.n1437 0.221854
R2782 VDPWR.n1362 VDPWR.n1361 0.221854
R2783 VDPWR.n1466 VDPWR.n1465 0.221854
R2784 VDPWR.n1346 VDPWR.n1345 0.221854
R2785 VDPWR.n1533 VDPWR 0.2005
R2786 VDPWR.n1392 VDPWR.n1387 0.199719
R2787 VDPWR.n126 VDPWR.n118 0.195812
R2788 VDPWR.n965 VDPWR.n964 0.189302
R2789 VDPWR.n960 VDPWR.n717 0.189302
R2790 VDPWR.n958 VDPWR.n957 0.189302
R2791 VDPWR.n953 VDPWR.n724 0.189302
R2792 VDPWR.n951 VDPWR.n950 0.189302
R2793 VDPWR.n946 VDPWR.n731 0.189302
R2794 VDPWR.n944 VDPWR.n943 0.189302
R2795 VDPWR.n939 VDPWR.n738 0.189302
R2796 VDPWR.n937 VDPWR.n936 0.189302
R2797 VDPWR.n932 VDPWR.n745 0.189302
R2798 VDPWR.n930 VDPWR.n929 0.189302
R2799 VDPWR.n925 VDPWR.n752 0.189302
R2800 VDPWR.n923 VDPWR.n922 0.189302
R2801 VDPWR.n918 VDPWR.n759 0.189302
R2802 VDPWR.n916 VDPWR.n915 0.189302
R2803 VDPWR.n911 VDPWR.n766 0.189302
R2804 VDPWR.n909 VDPWR.n908 0.189302
R2805 VDPWR.n904 VDPWR.n773 0.189302
R2806 VDPWR.n902 VDPWR.n901 0.189302
R2807 VDPWR.n897 VDPWR.n780 0.189302
R2808 VDPWR.n895 VDPWR.n894 0.189302
R2809 VDPWR.n890 VDPWR.n787 0.189302
R2810 VDPWR.n888 VDPWR.n887 0.189302
R2811 VDPWR.n883 VDPWR.n794 0.189302
R2812 VDPWR.n881 VDPWR.n880 0.189302
R2813 VDPWR.n876 VDPWR.n801 0.189302
R2814 VDPWR.n874 VDPWR.n873 0.189302
R2815 VDPWR.n869 VDPWR.n866 0.189302
R2816 VDPWR.n1564 VDPWR.n1563 0.189302
R2817 VDPWR.n1559 VDPWR.n1496 0.189302
R2818 VDPWR.n1557 VDPWR.n1556 0.189302
R2819 VDPWR.n1552 VDPWR.n1503 0.189302
R2820 VDPWR.n1550 VDPWR.n1549 0.189302
R2821 VDPWR.n1545 VDPWR.n1510 0.189302
R2822 VDPWR.n343 VDPWR.n340 0.189302
R2823 VDPWR.n349 VDPWR.n304 0.189302
R2824 VDPWR.n377 VDPWR.n374 0.189302
R2825 VDPWR.n383 VDPWR.n280 0.189302
R2826 VDPWR.n403 VDPWR.n400 0.189302
R2827 VDPWR.n409 VDPWR.n256 0.189302
R2828 VDPWR.n429 VDPWR.n426 0.189302
R2829 VDPWR.n435 VDPWR.n232 0.189302
R2830 VDPWR.n455 VDPWR.n452 0.189302
R2831 VDPWR.n461 VDPWR.n208 0.189302
R2832 VDPWR.n481 VDPWR.n478 0.189302
R2833 VDPWR.n487 VDPWR.n184 0.189302
R2834 VDPWR.n82 VDPWR.n37 0.189302
R2835 VDPWR.n110 VDPWR.n107 0.189302
R2836 VDPWR.n116 VDPWR.n13 0.189302
R2837 VDPWR.n1393 VDPWR.n1392 0.185396
R2838 VDPWR VDPWR.n501 0.182792
R2839 VDPWR VDPWR.n512 0.182792
R2840 VDPWR.n92 VDPWR.n84 0.182792
R2841 VDPWR VDPWR.n138 0.182792
R2842 VDPWR VDPWR.n149 0.182792
R2843 VDPWR.n359 VDPWR.n351 0.178885
R2844 VDPWR.n1393 VDPWR.n1334 0.174979
R2845 VDPWR.n127 VDPWR.n126 0.174979
R2846 VDPWR.n492 VDPWR.n491 0.166299
R2847 VDPWR.n503 VDPWR.n502 0.166299
R2848 VDPWR.n129 VDPWR.n128 0.166299
R2849 VDPWR.n140 VDPWR.n139 0.166299
R2850 VDPWR.n1334 VDPWR 0.164562
R2851 VDPWR.n1543 VDPWR.n1511 0.158052
R2852 VDPWR.n1535 VDPWR.n1528 0.158052
R2853 VDPWR.n76 VDPWR.n73 0.158052
R2854 VDPWR VDPWR.n1489 0.151542
R2855 VDPWR.n341 VDPWR.n304 0.141125
R2856 VDPWR.n375 VDPWR.n280 0.141125
R2857 VDPWR.n401 VDPWR.n256 0.141125
R2858 VDPWR.n427 VDPWR.n232 0.141125
R2859 VDPWR.n453 VDPWR.n208 0.141125
R2860 VDPWR.n479 VDPWR.n184 0.141125
R2861 VDPWR.n74 VDPWR.n37 0.141125
R2862 VDPWR.n108 VDPWR.n13 0.141125
R2863 VDPWR VDPWR.n1575 0.133312
R2864 VDPWR.n717 VDPWR.n712 0.13201
R2865 VDPWR.n959 VDPWR.n958 0.13201
R2866 VDPWR.n724 VDPWR.n719 0.13201
R2867 VDPWR.n952 VDPWR.n951 0.13201
R2868 VDPWR.n731 VDPWR.n726 0.13201
R2869 VDPWR.n945 VDPWR.n944 0.13201
R2870 VDPWR.n738 VDPWR.n733 0.13201
R2871 VDPWR.n938 VDPWR.n937 0.13201
R2872 VDPWR.n745 VDPWR.n740 0.13201
R2873 VDPWR.n931 VDPWR.n930 0.13201
R2874 VDPWR.n752 VDPWR.n747 0.13201
R2875 VDPWR.n924 VDPWR.n923 0.13201
R2876 VDPWR.n759 VDPWR.n754 0.13201
R2877 VDPWR.n917 VDPWR.n916 0.13201
R2878 VDPWR.n766 VDPWR.n761 0.13201
R2879 VDPWR.n910 VDPWR.n909 0.13201
R2880 VDPWR.n773 VDPWR.n768 0.13201
R2881 VDPWR.n903 VDPWR.n902 0.13201
R2882 VDPWR.n780 VDPWR.n775 0.13201
R2883 VDPWR.n896 VDPWR.n895 0.13201
R2884 VDPWR.n787 VDPWR.n782 0.13201
R2885 VDPWR.n889 VDPWR.n888 0.13201
R2886 VDPWR.n794 VDPWR.n789 0.13201
R2887 VDPWR.n882 VDPWR.n881 0.13201
R2888 VDPWR.n801 VDPWR.n796 0.13201
R2889 VDPWR.n875 VDPWR.n874 0.13201
R2890 VDPWR.n866 VDPWR.n803 0.13201
R2891 VDPWR.n868 VDPWR.n867 0.13201
R2892 VDPWR.n1496 VDPWR.n1491 0.13201
R2893 VDPWR.n1558 VDPWR.n1557 0.13201
R2894 VDPWR.n1503 VDPWR.n1498 0.13201
R2895 VDPWR.n1551 VDPWR.n1550 0.13201
R2896 VDPWR.n1510 VDPWR.n1505 0.13201
R2897 VDPWR.n342 VDPWR.n341 0.13201
R2898 VDPWR.n351 VDPWR.n350 0.13201
R2899 VDPWR.n376 VDPWR.n375 0.13201
R2900 VDPWR.n385 VDPWR.n384 0.13201
R2901 VDPWR.n402 VDPWR.n401 0.13201
R2902 VDPWR.n411 VDPWR.n410 0.13201
R2903 VDPWR.n428 VDPWR.n427 0.13201
R2904 VDPWR.n437 VDPWR.n436 0.13201
R2905 VDPWR.n454 VDPWR.n453 0.13201
R2906 VDPWR.n463 VDPWR.n462 0.13201
R2907 VDPWR.n480 VDPWR.n479 0.13201
R2908 VDPWR.n489 VDPWR.n488 0.13201
R2909 VDPWR.n75 VDPWR.n74 0.13201
R2910 VDPWR.n84 VDPWR.n83 0.13201
R2911 VDPWR.n109 VDPWR.n108 0.13201
R2912 VDPWR.n118 VDPWR.n117 0.13201
R2913 VDPWR.n339 VDPWR.n338 0.130708
R2914 VDPWR.n373 VDPWR.n372 0.130708
R2915 VDPWR.n399 VDPWR.n398 0.130708
R2916 VDPWR.n425 VDPWR.n424 0.130708
R2917 VDPWR.n451 VDPWR.n450 0.130708
R2918 VDPWR.n477 VDPWR.n476 0.130708
R2919 VDPWR.n72 VDPWR.n71 0.130708
R2920 VDPWR.n106 VDPWR.n105 0.130708
R2921 VDPWR.n526 VDPWR.n168 0.129176
R2922 VDPWR.n500 VDPWR.n499 0.127236
R2923 VDPWR.n511 VDPWR.n510 0.127236
R2924 VDPWR.n137 VDPWR.n136 0.127236
R2925 VDPWR.n148 VDPWR.n147 0.127236
R2926 VDPWR.n1533 VDPWR 0.1255
R2927 VDPWR.n1012 VDPWR.n1011 0.124275
R2928 VDPWR.n1030 VDPWR.n1029 0.124275
R2929 VDPWR.n1048 VDPWR.n1047 0.124275
R2930 VDPWR.n1066 VDPWR.n1065 0.124275
R2931 VDPWR.n1084 VDPWR.n1083 0.124275
R2932 VDPWR.n1102 VDPWR.n1101 0.124275
R2933 VDPWR.n1120 VDPWR.n1119 0.124275
R2934 VDPWR.n1138 VDPWR.n1137 0.124275
R2935 VDPWR.n535 VDPWR.n534 0.124275
R2936 VDPWR.n327 VDPWR 0.124198
R2937 VDPWR.n361 VDPWR 0.124198
R2938 VDPWR.n387 VDPWR 0.124198
R2939 VDPWR.n413 VDPWR 0.124198
R2940 VDPWR.n439 VDPWR 0.124198
R2941 VDPWR.n465 VDPWR 0.124198
R2942 VDPWR.n60 VDPWR 0.124198
R2943 VDPWR.n94 VDPWR 0.124198
R2944 VDPWR.n1010 VDPWR.n997 0.121824
R2945 VDPWR.n1028 VDPWR.n993 0.121824
R2946 VDPWR.n1046 VDPWR.n989 0.121824
R2947 VDPWR.n1064 VDPWR.n985 0.121824
R2948 VDPWR.n1082 VDPWR.n981 0.121824
R2949 VDPWR.n1100 VDPWR.n977 0.121824
R2950 VDPWR.n1118 VDPWR.n973 0.121824
R2951 VDPWR.n1136 VDPWR.n969 0.121824
R2952 VDPWR.n491 VDPWR.n178 0.115083
R2953 VDPWR.n502 VDPWR.n172 0.115083
R2954 VDPWR.n128 VDPWR.n7 0.115083
R2955 VDPWR.n139 VDPWR.n1 0.115083
R2956 VDPWR VDPWR.n1014 0.113245
R2957 VDPWR VDPWR.n1032 0.113245
R2958 VDPWR VDPWR.n1050 0.113245
R2959 VDPWR VDPWR.n1068 0.113245
R2960 VDPWR VDPWR.n1086 0.113245
R2961 VDPWR VDPWR.n1104 0.113245
R2962 VDPWR VDPWR.n1122 0.113245
R2963 VDPWR VDPWR.n1140 0.113245
R2964 VDPWR.n534 VDPWR.n533 0.110794
R2965 VDPWR.n533 VDPWR.n168 0.105892
R2966 VDPWR VDPWR.n1333 0.104667
R2967 VDPWR VDPWR.n525 0.103441
R2968 VDPWR.n1544 VDPWR.n1543 0.10076
R2969 VDPWR.n501 VDPWR.n500 0.0899097
R2970 VDPWR.n512 VDPWR.n511 0.0899097
R2971 VDPWR.n138 VDPWR.n137 0.0899097
R2972 VDPWR.n149 VDPWR.n148 0.0899097
R2973 VDPWR.n166 VDPWR.n165 0.0826078
R2974 VDPWR.n165 VDPWR.n162 0.0777059
R2975 VDPWR.n1565 VDPWR.n1564 0.0734167
R2976 VDPWR.n1575 VDPWR.n162 0.0715784
R2977 VDPWR.n1534 VDPWR.n1533 0.0708125
R2978 VDPWR.n1528 VDPWR.n1527 0.0708125
R2979 VDPWR.n867 VDPWR 0.0708125
R2980 VDPWR VDPWR.n339 0.0695104
R2981 VDPWR.n360 VDPWR 0.0695104
R2982 VDPWR VDPWR.n373 0.0695104
R2983 VDPWR.n386 VDPWR 0.0695104
R2984 VDPWR VDPWR.n399 0.0695104
R2985 VDPWR.n412 VDPWR 0.0695104
R2986 VDPWR VDPWR.n425 0.0695104
R2987 VDPWR.n438 VDPWR 0.0695104
R2988 VDPWR VDPWR.n451 0.0695104
R2989 VDPWR.n464 VDPWR 0.0695104
R2990 VDPWR VDPWR.n477 0.0695104
R2991 VDPWR VDPWR.n72 0.0695104
R2992 VDPWR.n93 VDPWR 0.0695104
R2993 VDPWR VDPWR.n106 0.0695104
R2994 VDPWR.n1569 VDPWR.n166 0.0666765
R2995 VDPWR.n499 VDPWR.n178 0.0647361
R2996 VDPWR.n510 VDPWR.n172 0.0647361
R2997 VDPWR.n136 VDPWR.n7 0.0647361
R2998 VDPWR.n147 VDPWR.n1 0.0647361
R2999 VDPWR.n357 VDPWR 0.063
R3000 VDPWR.n124 VDPWR 0.063
R3001 VDPWR.n90 VDPWR 0.063
R3002 VDPWR.n964 VDPWR.n712 0.0577917
R3003 VDPWR.n960 VDPWR.n959 0.0577917
R3004 VDPWR.n957 VDPWR.n719 0.0577917
R3005 VDPWR.n953 VDPWR.n952 0.0577917
R3006 VDPWR.n950 VDPWR.n726 0.0577917
R3007 VDPWR.n946 VDPWR.n945 0.0577917
R3008 VDPWR.n943 VDPWR.n733 0.0577917
R3009 VDPWR.n939 VDPWR.n938 0.0577917
R3010 VDPWR.n936 VDPWR.n740 0.0577917
R3011 VDPWR.n932 VDPWR.n931 0.0577917
R3012 VDPWR.n929 VDPWR.n747 0.0577917
R3013 VDPWR.n925 VDPWR.n924 0.0577917
R3014 VDPWR.n922 VDPWR.n754 0.0577917
R3015 VDPWR.n918 VDPWR.n917 0.0577917
R3016 VDPWR.n915 VDPWR.n761 0.0577917
R3017 VDPWR.n911 VDPWR.n910 0.0577917
R3018 VDPWR.n908 VDPWR.n768 0.0577917
R3019 VDPWR.n904 VDPWR.n903 0.0577917
R3020 VDPWR.n901 VDPWR.n775 0.0577917
R3021 VDPWR.n897 VDPWR.n896 0.0577917
R3022 VDPWR.n894 VDPWR.n782 0.0577917
R3023 VDPWR.n890 VDPWR.n889 0.0577917
R3024 VDPWR.n887 VDPWR.n789 0.0577917
R3025 VDPWR.n883 VDPWR.n882 0.0577917
R3026 VDPWR.n880 VDPWR.n796 0.0577917
R3027 VDPWR.n876 VDPWR.n875 0.0577917
R3028 VDPWR.n873 VDPWR.n803 0.0577917
R3029 VDPWR.n869 VDPWR.n868 0.0577917
R3030 VDPWR.n1563 VDPWR.n1491 0.0577917
R3031 VDPWR.n1559 VDPWR.n1558 0.0577917
R3032 VDPWR.n1556 VDPWR.n1498 0.0577917
R3033 VDPWR.n1552 VDPWR.n1551 0.0577917
R3034 VDPWR.n1549 VDPWR.n1505 0.0577917
R3035 VDPWR.n1545 VDPWR.n1544 0.0577917
R3036 VDPWR.n522 VDPWR.n515 0.0577917
R3037 VDPWR.n343 VDPWR.n342 0.0577917
R3038 VDPWR.n350 VDPWR.n349 0.0577917
R3039 VDPWR.n377 VDPWR.n376 0.0577917
R3040 VDPWR.n384 VDPWR.n383 0.0577917
R3041 VDPWR.n403 VDPWR.n402 0.0577917
R3042 VDPWR.n410 VDPWR.n409 0.0577917
R3043 VDPWR.n429 VDPWR.n428 0.0577917
R3044 VDPWR.n436 VDPWR.n435 0.0577917
R3045 VDPWR.n455 VDPWR.n454 0.0577917
R3046 VDPWR.n462 VDPWR.n461 0.0577917
R3047 VDPWR.n481 VDPWR.n480 0.0577917
R3048 VDPWR.n488 VDPWR.n487 0.0577917
R3049 VDPWR.n159 VDPWR.n152 0.0577917
R3050 VDPWR.n76 VDPWR.n75 0.0577917
R3051 VDPWR.n83 VDPWR.n82 0.0577917
R3052 VDPWR.n110 VDPWR.n109 0.0577917
R3053 VDPWR.n117 VDPWR.n116 0.0577917
R3054 VDPWR.n513 VDPWR 0.0439028
R3055 VDPWR.n150 VDPWR 0.0439028
R3056 VDPWR.n591 VDPWR.n574 0.0432215
R3057 VDPWR.n608 VDPWR.n569 0.0432215
R3058 VDPWR.n625 VDPWR.n564 0.0432215
R3059 VDPWR.n642 VDPWR.n559 0.0432215
R3060 VDPWR.n659 VDPWR.n554 0.0432215
R3061 VDPWR.n676 VDPWR.n549 0.0432215
R3062 VDPWR.n693 VDPWR.n544 0.0432215
R3063 VDPWR.n710 VDPWR.n539 0.0432215
R3064 VDPWR VDPWR.n490 0.0421667
R3065 VDPWR VDPWR.n127 0.0421667
R3066 VDPWR.n170 VDPWR 0.0295179
R3067 VDPWR.n1527 VDPWR.n1511 0.0278438
R3068 VDPWR.n1535 VDPWR.n1534 0.0278438
R3069 VDPWR.n1575 VDPWR 0.0201078
R3070 VDPWR.n1333 VDPWR 0.0187292
R3071 VDPWR.n526 VDPWR 0.0103039
R3072 VDPWR VDPWR.n360 0.00701042
R3073 VDPWR VDPWR.n386 0.00701042
R3074 VDPWR VDPWR.n412 0.00701042
R3075 VDPWR VDPWR.n438 0.00701042
R3076 VDPWR VDPWR.n464 0.00701042
R3077 VDPWR VDPWR.n93 0.00701042
R3078 VDPWR.n523 VDPWR.n522 0.00440625
R3079 VDPWR.n160 VDPWR.n159 0.00440625
R3080 VDPWR.n1011 VDPWR.n1010 0.00295098
R3081 VDPWR.n1029 VDPWR.n1028 0.00295098
R3082 VDPWR.n1047 VDPWR.n1046 0.00295098
R3083 VDPWR.n1065 VDPWR.n1064 0.00295098
R3084 VDPWR.n1083 VDPWR.n1082 0.00295098
R3085 VDPWR.n1101 VDPWR.n1100 0.00295098
R3086 VDPWR.n1119 VDPWR.n1118 0.00295098
R3087 VDPWR.n1137 VDPWR.n1136 0.00295098
R3088 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 784.053
R3089 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 784.053
R3090 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 784.053
R3091 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 784.053
R3092 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 539.841
R3093 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 539.841
R3094 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 539.841
R3095 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 539.841
R3096 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 215.293
R3097 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 215.293
R3098 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 215.293
R3099 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 215.293
R3100 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 168.659
R3101 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 167.992
R3102 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 166.144
R3103 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 165.8
R3104 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 85.2499
R3105 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 85.2499
R3106 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 83.7172
R3107 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 83.7172
R3108 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 75.7282
R3109 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 66.3172
R3110 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 36.1505
R3111 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 36.1505
R3112 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 34.5438
R3113 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 34.5438
R3114 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 17.4005
R3115 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 17.4005
R3116 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 17.2391
R3117 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 9.52217
R3118 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 9.52217
R3119 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 6.39571
R3120 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 5.30824
R3121 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 4.94887
R3122 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 1.48097
R3123 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 1.06691
R3124 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.539562
R3125 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.391125
R3126 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 0.160656
R3127 tdc_0.start_buffer_0.start_buff.n11 tdc_0.start_buffer_0.start_buff.t21 543.053
R3128 tdc_0.start_buffer_0.start_buff.n12 tdc_0.start_buffer_0.start_buff.t16 543.053
R3129 tdc_0.start_buffer_0.start_buff.n10 tdc_0.start_buffer_0.start_buff.t10 543.053
R3130 tdc_0.start_buffer_0.start_buff.n1 tdc_0.start_buffer_0.start_buff.t11 539.841
R3131 tdc_0.start_buffer_0.start_buff.n0 tdc_0.start_buffer_0.start_buff.t15 539.841
R3132 tdc_0.start_buffer_0.start_buff.n4 tdc_0.start_buffer_0.start_buff.t13 539.841
R3133 tdc_0.start_buffer_0.start_buff.n3 tdc_0.start_buffer_0.start_buff.t19 539.841
R3134 tdc_0.start_buffer_0.start_buff.n11 tdc_0.start_buffer_0.start_buff.t18 221.72
R3135 tdc_0.start_buffer_0.start_buff.n12 tdc_0.start_buffer_0.start_buff.t14 221.72
R3136 tdc_0.start_buffer_0.start_buff.n10 tdc_0.start_buffer_0.start_buff.t22 221.72
R3137 tdc_0.start_buffer_0.start_buff.n13 tdc_0.start_buffer_0.start_buff.n11 218.32
R3138 tdc_0.start_buffer_0.start_buff.n13 tdc_0.start_buffer_0.start_buff.n12 217.734
R3139 tdc_0.start_buffer_0.start_buff.n1 tdc_0.start_buffer_0.start_buff.t20 215.293
R3140 tdc_0.start_buffer_0.start_buff.n0 tdc_0.start_buffer_0.start_buff.t12 215.293
R3141 tdc_0.start_buffer_0.start_buff.n4 tdc_0.start_buffer_0.start_buff.t23 215.293
R3142 tdc_0.start_buffer_0.start_buff.n3 tdc_0.start_buffer_0.start_buff.t17 215.293
R3143 tdc_0.start_buffer_0.start_buff.n14 tdc_0.start_buffer_0.start_buff.n10 213.234
R3144 tdc_0.start_buffer_0.start_buff.n6 tdc_0.start_buffer_0.start_buff.n2 166.149
R3145 tdc_0.start_buffer_0.start_buff.n6 tdc_0.start_buffer_0.start_buff.n5 165.8
R3146 tdc_0.start_buffer_0.start_buff.n18 tdc_0.start_buffer_0.start_buff.t4 85.2499
R3147 tdc_0.start_buffer_0.start_buff.n17 tdc_0.start_buffer_0.start_buff.t6 85.2499
R3148 tdc_0.start_buffer_0.start_buff.n20 tdc_0.start_buffer_0.start_buff.t7 85.2499
R3149 tdc_0.start_buffer_0.start_buff.n7 tdc_0.start_buffer_0.start_buff.t9 85.1574
R3150 tdc_0.start_buffer_0.start_buff.n9 tdc_0.start_buffer_0.start_buff.t5 83.8097
R3151 tdc_0.start_buffer_0.start_buff.n7 tdc_0.start_buffer_0.start_buff.t8 83.8097
R3152 tdc_0.start_buffer_0.start_buff.n20 tdc_0.start_buffer_0.start_buff.t3 83.7172
R3153 tdc_0.start_buffer_0.start_buff.n16 tdc_0.start_buffer_0.start_buff.t1 83.7172
R3154 tdc_0.start_buffer_0.start_buff.n18 tdc_0.start_buffer_0.start_buff.t0 83.7172
R3155 tdc_0.start_buffer_0.start_buff.n17 tdc_0.start_buffer_0.start_buff.t2 83.7172
R3156 tdc_0.start_buffer_0.start_buff.n2 tdc_0.start_buffer_0.start_buff.n1 36.1505
R3157 tdc_0.start_buffer_0.start_buff.n5 tdc_0.start_buffer_0.start_buff.n3 36.1505
R3158 tdc_0.start_buffer_0.start_buff.n2 tdc_0.start_buffer_0.start_buff.n0 34.5438
R3159 tdc_0.start_buffer_0.start_buff.n5 tdc_0.start_buffer_0.start_buff.n4 34.5438
R3160 tdc_0.start_buffer_0.start_buff.n8 tdc_0.start_buffer_0.start_buff.n6 11.8364
R3161 tdc_0.start_buffer_0.start_buff.n9 tdc_0.start_buffer_0.start_buff 8.40722
R3162 tdc_0.start_buffer_0.start_buff.n8 tdc_0.start_buffer_0.start_buff.n7 5.74235
R3163 tdc_0.start_buffer_0.start_buff.n19 tdc_0.start_buffer_0.start_buff.n17 5.16238
R3164 tdc_0.start_buffer_0.start_buff.n14 tdc_0.start_buffer_0.start_buff.n13 5.08518
R3165 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_buff.n16 4.70702
R3166 tdc_0.start_buffer_0.start_buff.n19 tdc_0.start_buffer_0.start_buff.n18 4.64452
R3167 tdc_0.start_buffer_0.start_buff.n21 tdc_0.start_buffer_0.start_buff.n20 4.64452
R3168 tdc_0.start_buffer_0.start_buff.n15 tdc_0.start_buffer_0.start_buff.n9 0.918978
R3169 tdc_0.start_buffer_0.start_buff.n21 tdc_0.start_buffer_0.start_buff.n19 0.518357
R3170 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_buff.n21 0.455857
R3171 tdc_0.start_buffer_0.start_buff.n16 tdc_0.start_buffer_0.start_buff.n15 0.3755
R3172 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_buff.n8 0.285656
R3173 tdc_0.start_buffer_0.start_buff.n15 tdc_0.start_buffer_0.start_buff.n14 0.247513
R3174 tdc_0.start_buffer_0.start_delay.n1 tdc_0.start_buffer_0.start_delay.t14 539.841
R3175 tdc_0.start_buffer_0.start_delay.n0 tdc_0.start_buffer_0.start_delay.t8 539.841
R3176 tdc_0.start_buffer_0.start_delay.n4 tdc_0.start_buffer_0.start_delay.t10 539.841
R3177 tdc_0.start_buffer_0.start_delay.n3 tdc_0.start_buffer_0.start_delay.t13 539.841
R3178 tdc_0.start_buffer_0.start_delay.n1 tdc_0.start_buffer_0.start_delay.t12 215.293
R3179 tdc_0.start_buffer_0.start_delay.n0 tdc_0.start_buffer_0.start_delay.t15 215.293
R3180 tdc_0.start_buffer_0.start_delay.n4 tdc_0.start_buffer_0.start_delay.t9 215.293
R3181 tdc_0.start_buffer_0.start_delay.n3 tdc_0.start_buffer_0.start_delay.t11 215.293
R3182 tdc_0.start_buffer_0.start_delay.n6 tdc_0.start_buffer_0.start_delay.n2 166.144
R3183 tdc_0.start_buffer_0.start_delay.n6 tdc_0.start_buffer_0.start_delay.n5 165.8
R3184 tdc_0.start_buffer_0.start_delay.n9 tdc_0.start_buffer_0.start_delay.t4 85.2499
R3185 tdc_0.start_buffer_0.start_delay.n7 tdc_0.start_buffer_0.start_delay.t5 85.2499
R3186 tdc_0.start_buffer_0.start_delay.n8 tdc_0.start_buffer_0.start_delay.t6 85.2499
R3187 tdc_0.start_buffer_0.start_delay.n11 tdc_0.start_buffer_0.start_delay.t3 84.7281
R3188 tdc_0.start_buffer_0.start_delay.n8 tdc_0.start_buffer_0.start_delay.t1 83.7172
R3189 tdc_0.start_buffer_0.start_delay.n12 tdc_0.start_buffer_0.start_delay.t2 83.7172
R3190 tdc_0.start_buffer_0.start_delay.n9 tdc_0.start_buffer_0.start_delay.t7 83.7172
R3191 tdc_0.start_buffer_0.start_delay.n7 tdc_0.start_buffer_0.start_delay.t0 83.7172
R3192 tdc_0.start_buffer_0.start_delay.n2 tdc_0.start_buffer_0.start_delay.n0 36.1505
R3193 tdc_0.start_buffer_0.start_delay.n5 tdc_0.start_buffer_0.start_delay.n3 36.1505
R3194 tdc_0.start_buffer_0.start_delay.n2 tdc_0.start_buffer_0.start_delay.n1 34.5438
R3195 tdc_0.start_buffer_0.start_delay.n5 tdc_0.start_buffer_0.start_delay.n4 34.5438
R3196 tdc_0.start_buffer_0.start_delay tdc_0.start_buffer_0.start_delay.n7 6.45821
R3197 tdc_0.start_buffer_0.start_delay.n10 tdc_0.start_buffer_0.start_delay.n8 5.16238
R3198 tdc_0.start_buffer_0.start_delay.n13 tdc_0.start_buffer_0.start_delay.n12 4.64452
R3199 tdc_0.start_buffer_0.start_delay.n10 tdc_0.start_buffer_0.start_delay.n9 4.64452
R3200 tdc_0.start_buffer_0.start_delay.n14 tdc_0.start_buffer_0.start_delay.n13 0.759429
R3201 tdc_0.start_buffer_0.start_delay.n13 tdc_0.start_buffer_0.start_delay.n10 0.518357
R3202 tdc_0.start_buffer_0.start_delay.n14 tdc_0.start_buffer_0.start_delay 0.471203
R3203 tdc_0.start_buffer_0.start_delay tdc_0.start_buffer_0.start_delay.n6 0.46925
R3204 tdc_0.start_buffer_0.start_delay.n12 tdc_0.start_buffer_0.start_delay.n11 0.3755
R3205 tdc_0.start_buffer_0.start_delay.n11 tdc_0.start_buffer_0.start_delay 0.234296
R3206 tdc_0.start_buffer_0.start_delay tdc_0.start_buffer_0.start_delay.n14 0.127453
R3207 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t2 628.097
R3208 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t6 622.766
R3209 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t4 523.774
R3210 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t5 304.647
R3211 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t7 304.647
R3212 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t3 202.44
R3213 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 169.062
R3214 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 166.237
R3215 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t0 84.7557
R3216 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t1 84.1197
R3217 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 12.6535
R3218 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 5.48979
R3219 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en 4.5005
R3220 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 1.09595
R3221 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 890.727
R3222 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 742.783
R3223 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 641.061
R3224 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 623.388
R3225 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 547.874
R3226 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 431.807
R3227 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 427.875
R3228 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 340.632
R3229 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 208.631
R3230 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 168.007
R3231 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R3232 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 31.2103
R3233 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 31.0962
R3234 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 9.52217
R3235 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R3236 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 8.91506
R3237 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R3238 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R3239 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R3240 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R3241 VGND.n1747 VGND.n166 145435
R3242 VGND.n1747 VGND.n1746 89027.6
R3243 VGND.n316 VGND.n188 35396
R3244 VGND.n1004 VGND.n166 35396
R3245 VGND.n1747 VGND.n167 31825.6
R3246 VGND.n146 VGND.n135 24188.9
R3247 VGND.n315 VGND.n137 22872.1
R3248 VGND.n1828 VGND.t0 18604.5
R3249 VGND.n168 VGND.n167 16815
R3250 VGND.n208 VGND.n188 16612
R3251 VGND.n1712 VGND.n331 14632.6
R3252 VGND.n208 VGND.t0 14477.4
R3253 VGND.n1577 VGND.t259 13628.8
R3254 VGND.n1826 VGND.t0 11061.3
R3255 VGND.n1569 VGND.n1568 9459.64
R3256 VGND.n330 VGND.n167 9082.84
R3257 VGND.n1761 VGND.t8 7799.94
R3258 VGND.n1794 VGND.n5 6289.43
R3259 VGND.n1578 VGND.n1577 6212.87
R3260 VGND.n1828 VGND.n1827 5291.8
R3261 VGND.n1577 VGND.n5 4980.04
R3262 VGND.n1709 VGND.n1578 4836.21
R3263 VGND.t236 VGND.n1828 4811.74
R3264 VGND.n314 VGND.n189 4594.02
R3265 VGND.n1569 VGND.n563 4479.04
R3266 VGND.n1570 VGND.n562 4479.04
R3267 VGND.n1571 VGND.n561 4479.04
R3268 VGND.n1572 VGND.n560 4479.04
R3269 VGND.n1573 VGND.n559 4479.04
R3270 VGND.n1574 VGND.n558 4479.04
R3271 VGND.n1575 VGND.n557 4479.04
R3272 VGND.n1576 VGND.n556 4479.04
R3273 VGND.n857 VGND.n138 4447.27
R3274 VGND.n1760 VGND.n139 4447.27
R3275 VGND.n260 VGND.n259 4447.27
R3276 VGND.n227 VGND.n226 4447.27
R3277 VGND.n1034 VGND.n520 4283.98
R3278 VGND.n1018 VGND.n520 4283.98
R3279 VGND.n696 VGND.n520 4283.98
R3280 VGND.n678 VGND.n520 4283.98
R3281 VGND.n654 VGND.n520 4283.98
R3282 VGND.n630 VGND.n520 4283.98
R3283 VGND.n606 VGND.n520 4283.98
R3284 VGND.t234 VGND.n1761 4154.59
R3285 VGND.n1548 VGND.n1163 3781.58
R3286 VGND.n1548 VGND.n1164 3781.58
R3287 VGND.n1548 VGND.n1165 3781.58
R3288 VGND.n1548 VGND.n1166 3781.58
R3289 VGND.n1548 VGND.n1167 3781.58
R3290 VGND.n1549 VGND.n1548 3781.58
R3291 VGND.n1548 VGND.n1547 3781.58
R3292 VGND.n1746 VGND.n331 3732.45
R3293 VGND.n1749 VGND.n138 3442.57
R3294 VGND.n1760 VGND.n140 3442.57
R3295 VGND.n259 VGND.n256 3442.57
R3296 VGND.n254 VGND.n227 3442.57
R3297 VGND.n1147 VGND.n563 3439.59
R3298 VGND.n331 VGND.n6 3358.06
R3299 VGND.n857 VGND.n161 3165.68
R3300 VGND.n157 VGND.n139 3165.68
R3301 VGND.n260 VGND.n220 3165.68
R3302 VGND.n230 VGND.n226 3165.68
R3303 VGND.n1161 VGND.n563 3093.4
R3304 VGND.n1470 VGND.n562 3093.4
R3305 VGND.n1458 VGND.n561 3093.4
R3306 VGND.n1446 VGND.n560 3093.4
R3307 VGND.n1434 VGND.n559 3093.4
R3308 VGND.n1422 VGND.n558 3093.4
R3309 VGND.n1409 VGND.n557 3093.4
R3310 VGND.n1535 VGND.n556 3093.4
R3311 VGND.n1236 VGND.n521 3089.56
R3312 VGND.n1386 VGND.n527 3089.56
R3313 VGND.n1376 VGND.n522 3089.56
R3314 VGND.n1351 VGND.n526 3089.56
R3315 VGND.n1326 VGND.n523 3089.56
R3316 VGND.n1301 VGND.n525 3089.56
R3317 VGND.n1727 VGND.n519 3089.56
R3318 VGND.n1725 VGND.n529 3089.56
R3319 VGND.n1235 VGND.n1170 2843.1
R3320 VGND.n1385 VGND.n1171 2843.1
R3321 VGND.n1375 VGND.n1172 2843.1
R3322 VGND.n1350 VGND.n1173 2843.1
R3323 VGND.n1325 VGND.n1174 2843.1
R3324 VGND.n1300 VGND.n1175 2843.1
R3325 VGND.n1177 VGND.n1176 2843.1
R3326 VGND.n1169 VGND.n536 2843.1
R3327 VGND.n1827 VGND.n1826 2773.54
R3328 VGND.n1711 VGND.n1710 2755.48
R3329 VGND.n1568 VGND.n565 2713.47
R3330 VGND.n314 VGND.n313 2502.61
R3331 VGND.n331 VGND.n330 2480.88
R3332 VGND.n1568 VGND.n1567 2378.68
R3333 VGND.n1240 VGND.n521 2350.81
R3334 VGND.n1226 VGND.n527 2350.81
R3335 VGND.n1365 VGND.n522 2350.81
R3336 VGND.n1340 VGND.n526 2350.81
R3337 VGND.n1315 VGND.n523 2350.81
R3338 VGND.n1290 VGND.n525 2350.81
R3339 VGND.n1727 VGND.n518 2350.81
R3340 VGND.n1725 VGND.n528 2350.81
R3341 VGND.n1749 VGND.n162 2206.4
R3342 VGND.n158 VGND.n140 2206.4
R3343 VGND.n256 VGND.n223 2206.4
R3344 VGND.n254 VGND.n225 2206.4
R3345 VGND.n238 VGND.n136 2152.16
R3346 VGND.n151 VGND.n146 2067.34
R3347 VGND.n1600 VGND.n1595 2058.56
R3348 VGND.n1693 VGND.n1595 2058.56
R3349 VGND.n1690 VGND.n1603 2058.56
R3350 VGND.n1622 VGND.n1603 2058.56
R3351 VGND.n1624 VGND.n1619 2058.56
R3352 VGND.n1675 VGND.n1619 2058.56
R3353 VGND.n1672 VGND.n1627 2058.56
R3354 VGND.n1649 VGND.n1627 2058.56
R3355 VGND.n1651 VGND.n1646 2058.56
R3356 VGND.n1657 VGND.n1646 2058.56
R3357 VGND.n1792 VGND.n75 2058.56
R3358 VGND.n1654 VGND.n75 2058.56
R3359 VGND.n1598 VGND.n1579 2058.56
R3360 VGND.n1707 VGND.n1579 2058.56
R3361 VGND.n1566 VGND.n566 2058.56
R3362 VGND.n1148 VGND.n566 2058.56
R3363 VGND.n1160 VGND.n1159 2058.56
R3364 VGND.n1551 VGND.n1159 2058.56
R3365 VGND.n1471 VGND.n1466 2058.56
R3366 VGND.n1467 VGND.n1466 2058.56
R3367 VGND.n1459 VGND.n1454 2058.56
R3368 VGND.n1455 VGND.n1454 2058.56
R3369 VGND.n1447 VGND.n1442 2058.56
R3370 VGND.n1443 VGND.n1442 2058.56
R3371 VGND.n1435 VGND.n1430 2058.56
R3372 VGND.n1431 VGND.n1430 2058.56
R3373 VGND.n1423 VGND.n1418 2058.56
R3374 VGND.n1419 VGND.n1418 2058.56
R3375 VGND.n1410 VGND.n1401 2058.56
R3376 VGND.n1545 VGND.n1401 2058.56
R3377 VGND.n1533 VGND.n1532 2058.56
R3378 VGND.n1534 VGND.n1533 2058.56
R3379 VGND.n1189 VGND.n1188 2029.1
R3380 VGND.n1393 VGND.n1220 2029.1
R3381 VGND.n1192 VGND.n1191 2029.1
R3382 VGND.n1218 VGND.n1217 2029.1
R3383 VGND.n1195 VGND.n1194 2029.1
R3384 VGND.n1215 VGND.n1214 2029.1
R3385 VGND.n1212 VGND.n1197 2029.1
R3386 VGND.n1395 VGND.n1186 2029.1
R3387 VGND.n1251 VGND.n1184 1929.2
R3388 VGND.n1230 VGND.n1183 1929.2
R3389 VGND.n1366 VGND.n1182 1929.2
R3390 VGND.n1341 VGND.n1181 1929.2
R3391 VGND.n1316 VGND.n1180 1929.2
R3392 VGND.n1291 VGND.n1179 1929.2
R3393 VGND.n1204 VGND.n1178 1929.2
R3394 VGND.n1399 VGND.n1185 1929.2
R3395 VGND.n509 VGND.n6 1814.76
R3396 VGND.n1549 VGND.n562 1809.14
R3397 VGND.n1167 VGND.n561 1809.14
R3398 VGND.n1166 VGND.n560 1809.14
R3399 VGND.n1165 VGND.n559 1809.14
R3400 VGND.n1164 VGND.n558 1809.14
R3401 VGND.n1163 VGND.n557 1809.14
R3402 VGND.n1547 VGND.n556 1809.14
R3403 VGND.n1568 VGND.n564 1741.86
R3404 VGND.n1189 VGND.n1187 1718.82
R3405 VGND.n1393 VGND.n1219 1718.82
R3406 VGND.n1192 VGND.n1190 1718.82
R3407 VGND.n1218 VGND.n1216 1718.82
R3408 VGND.n1195 VGND.n1193 1718.82
R3409 VGND.n1215 VGND.n1213 1718.82
R3410 VGND.n1212 VGND.n1196 1718.82
R3411 VGND.n1395 VGND.n535 1718.82
R3412 VGND.n1763 VGND.n135 1708.68
R3413 VGND.n1829 VGND.n3 1707.33
R3414 VGND.n1831 VGND.n3 1707.33
R3415 VGND.n1764 VGND.n133 1707.33
R3416 VGND.n1764 VGND.n134 1707.33
R3417 VGND.n188 VGND.n6 1644.04
R3418 VGND.n1550 VGND.n1549 1630.46
R3419 VGND.n1468 VGND.n1167 1630.46
R3420 VGND.n1456 VGND.n1166 1630.46
R3421 VGND.n1444 VGND.n1165 1630.46
R3422 VGND.n1432 VGND.n1164 1630.46
R3423 VGND.n1420 VGND.n1163 1630.46
R3424 VGND.n1547 VGND.n1546 1630.46
R3425 VGND.n185 VGND.n180 1626.7
R3426 VGND.n318 VGND.n180 1626.7
R3427 VGND.n312 VGND.n192 1626.7
R3428 VGND.n312 VGND.n193 1626.7
R3429 VGND.n302 VGND.n190 1626.7
R3430 VGND.n304 VGND.n190 1626.7
R3431 VGND.n1000 VGND.n737 1626.7
R3432 VGND.n1006 VGND.n737 1626.7
R3433 VGND.n975 VGND.n770 1626.7
R3434 VGND.n977 VGND.n770 1626.7
R3435 VGND.n974 VGND.n790 1626.7
R3436 VGND.n790 VGND.n772 1626.7
R3437 VGND.n953 VGND.n789 1626.7
R3438 VGND.n953 VGND.n773 1626.7
R3439 VGND.n808 VGND.n788 1626.7
R3440 VGND.n808 VGND.n774 1626.7
R3441 VGND.n931 VGND.n787 1626.7
R3442 VGND.n931 VGND.n775 1626.7
R3443 VGND.n822 VGND.n786 1626.7
R3444 VGND.n822 VGND.n776 1626.7
R3445 VGND.n909 VGND.n785 1626.7
R3446 VGND.n909 VGND.n777 1626.7
R3447 VGND.n836 VGND.n784 1626.7
R3448 VGND.n836 VGND.n778 1626.7
R3449 VGND.n887 VGND.n783 1626.7
R3450 VGND.n887 VGND.n779 1626.7
R3451 VGND.n850 VGND.n782 1626.7
R3452 VGND.n850 VGND.n780 1626.7
R3453 VGND.n1016 VGND.n726 1626.7
R3454 VGND.n998 VGND.n726 1626.7
R3455 VGND.n328 VGND.n169 1626.7
R3456 VGND.n183 VGND.n169 1626.7
R3457 VGND.n1761 VGND.n136 1617.44
R3458 VGND.n1253 VGND.n1240 1562.99
R3459 VGND.n1232 VGND.n1226 1562.99
R3460 VGND.n1368 VGND.n1365 1562.99
R3461 VGND.n1343 VGND.n1340 1562.99
R3462 VGND.n1318 VGND.n1315 1562.99
R3463 VGND.n1293 VGND.n1290 1562.99
R3464 VGND.n1202 VGND.n518 1562.99
R3465 VGND.n1714 VGND.n528 1562.99
R3466 VGND.n1570 VGND.n1569 1482.26
R3467 VGND.n1571 VGND.n1570 1482.26
R3468 VGND.n1572 VGND.n1571 1482.26
R3469 VGND.n1573 VGND.n1572 1482.26
R3470 VGND.n1574 VGND.n1573 1482.26
R3471 VGND.n1575 VGND.n1574 1482.26
R3472 VGND.n1576 VGND.n1575 1482.26
R3473 VGND.n1578 VGND.n1576 1458.22
R3474 VGND.n1753 VGND.n162 1438.1
R3475 VGND.n1755 VGND.n158 1438.1
R3476 VGND.n264 VGND.n223 1438.1
R3477 VGND.n225 VGND.n224 1438.1
R3478 VGND.n1793 VGND.n1791 1396.01
R3479 VGND.n1825 VGND.n1824 1325.13
R3480 VGND.n1710 VGND.n555 1263.93
R3481 VGND.n1709 VGND.n1708 1228.29
R3482 VGND.n1188 VGND.n1184 1210.97
R3483 VGND.n1220 VGND.n1183 1210.97
R3484 VGND.n1191 VGND.n1182 1210.97
R3485 VGND.n1217 VGND.n1181 1210.97
R3486 VGND.n1194 VGND.n1180 1210.97
R3487 VGND.n1214 VGND.n1179 1210.97
R3488 VGND.n1197 VGND.n1178 1210.97
R3489 VGND.n1399 VGND.n1186 1210.97
R3490 VGND.n1188 VGND.n1170 1199.38
R3491 VGND.n1220 VGND.n1171 1199.38
R3492 VGND.n1191 VGND.n1172 1199.38
R3493 VGND.n1217 VGND.n1173 1199.38
R3494 VGND.n1194 VGND.n1174 1199.38
R3495 VGND.n1214 VGND.n1175 1199.38
R3496 VGND.n1197 VGND.n1177 1199.38
R3497 VGND.n1186 VGND.n1169 1199.38
R3498 VGND.n1827 VGND.n5 1074.72
R3499 VGND.n1753 VGND.n161 1065.44
R3500 VGND.n1755 VGND.n157 1065.44
R3501 VGND.n264 VGND.n220 1065.44
R3502 VGND.n230 VGND.n224 1065.44
R3503 VGND.n300 VGND.n283 1058.19
R3504 VGND.n283 VGND.n204 1058.19
R3505 VGND.n288 VGND.n282 1058.19
R3506 VGND.n288 VGND.n205 1058.19
R3507 VGND.n281 VGND.n210 1058.19
R3508 VGND.n210 VGND.n206 1058.19
R3509 VGND.n215 VGND.n209 1058.19
R3510 VGND.n215 VGND.n207 1058.19
R3511 VGND.n240 VGND.n237 1058.19
R3512 VGND.n242 VGND.n237 1058.19
R3513 VGND.n152 VGND.n145 1058.19
R3514 VGND.n150 VGND.n145 1058.19
R3515 VGND.n989 VGND.n740 1058.19
R3516 VGND.n991 VGND.n740 1058.19
R3517 VGND.n988 VGND.n763 1058.19
R3518 VGND.n763 VGND.n742 1058.19
R3519 VGND.n797 VGND.n762 1058.19
R3520 VGND.n797 VGND.n743 1058.19
R3521 VGND.n800 VGND.n761 1058.19
R3522 VGND.n800 VGND.n744 1058.19
R3523 VGND.n811 VGND.n760 1058.19
R3524 VGND.n811 VGND.n745 1058.19
R3525 VGND.n814 VGND.n759 1058.19
R3526 VGND.n814 VGND.n746 1058.19
R3527 VGND.n825 VGND.n758 1058.19
R3528 VGND.n825 VGND.n747 1058.19
R3529 VGND.n828 VGND.n757 1058.19
R3530 VGND.n828 VGND.n748 1058.19
R3531 VGND.n839 VGND.n756 1058.19
R3532 VGND.n839 VGND.n749 1058.19
R3533 VGND.n842 VGND.n755 1058.19
R3534 VGND.n842 VGND.n750 1058.19
R3535 VGND.n853 VGND.n754 1058.19
R3536 VGND.n853 VGND.n751 1058.19
R3537 VGND.n856 VGND.n753 1058.19
R3538 VGND.n856 VGND.n752 1058.19
R3539 VGND.n1804 VGND.n12 1058.19
R3540 VGND.n510 VGND.n343 1058.19
R3541 VGND.n1773 VGND.n79 1058.19
R3542 VGND.n1790 VGND.n84 1058.19
R3543 VGND.n1826 VGND.n1825 987.279
R3544 VGND.n1567 VGND.t146 815.229
R3545 VGND.n1146 VGND.t457 815.229
R3546 VGND.t417 VGND.n1146 815.229
R3547 VGND.n1147 VGND.t419 815.229
R3548 VGND.t333 VGND.n1161 815.229
R3549 VGND.n1162 VGND.t498 815.229
R3550 VGND.t209 VGND.n1162 815.229
R3551 VGND.n1550 VGND.t75 815.229
R3552 VGND.n1470 VGND.t350 815.229
R3553 VGND.t352 VGND.n1469 815.229
R3554 VGND.n1469 VGND.t340 815.229
R3555 VGND.t338 VGND.n1468 815.229
R3556 VGND.n1458 VGND.t519 815.229
R3557 VGND.t136 VGND.n1457 815.229
R3558 VGND.n1457 VGND.t69 815.229
R3559 VGND.t104 VGND.n1456 815.229
R3560 VGND.n1446 VGND.t447 815.229
R3561 VGND.t152 VGND.n1445 815.229
R3562 VGND.n1445 VGND.t388 815.229
R3563 VGND.t386 VGND.n1444 815.229
R3564 VGND.n1434 VGND.t408 815.229
R3565 VGND.t414 VGND.n1433 815.229
R3566 VGND.n1433 VGND.t272 815.229
R3567 VGND.t312 VGND.n1432 815.229
R3568 VGND.n1422 VGND.t310 815.229
R3569 VGND.t52 VGND.n1421 815.229
R3570 VGND.n1421 VGND.t17 815.229
R3571 VGND.t19 VGND.n1420 815.229
R3572 VGND.n1409 VGND.t556 815.229
R3573 VGND.t119 VGND.n1408 815.229
R3574 VGND.n1408 VGND.t440 815.229
R3575 VGND.n1546 VGND.t211 815.229
R3576 VGND.t65 VGND.n1535 815.229
R3577 VGND.n1536 VGND.t79 815.229
R3578 VGND.n1536 VGND.t102 815.229
R3579 VGND.n62 VGND.n61 760.639
R3580 VGND.n56 VGND.n55 760.639
R3581 VGND.n50 VGND.n49 760.639
R3582 VGND.n44 VGND.n43 760.639
R3583 VGND.n38 VGND.n37 760.639
R3584 VGND.n32 VGND.n31 760.639
R3585 VGND.n26 VGND.n25 760.639
R3586 VGND.n470 VGND.n16 760.639
R3587 VGND.n466 VGND.n465 760.639
R3588 VGND.n460 VGND.n459 760.639
R3589 VGND.n454 VGND.n453 760.639
R3590 VGND.n448 VGND.n447 760.639
R3591 VGND.n442 VGND.n441 760.639
R3592 VGND.n436 VGND.n435 760.639
R3593 VGND.n430 VGND.n429 760.639
R3594 VGND.n424 VGND.n423 760.639
R3595 VGND.n418 VGND.n417 760.639
R3596 VGND.n412 VGND.n411 760.639
R3597 VGND.n406 VGND.n405 760.639
R3598 VGND.n400 VGND.n399 760.639
R3599 VGND.n394 VGND.n393 760.639
R3600 VGND.n388 VGND.n387 760.639
R3601 VGND.n382 VGND.n381 760.639
R3602 VGND.n376 VGND.n364 760.639
R3603 VGND.n366 VGND.n363 760.639
R3604 VGND.n368 VGND.n344 760.639
R3605 VGND.n20 VGND.n17 760.639
R3606 VGND.n124 VGND.n123 760.639
R3607 VGND.n118 VGND.n117 760.639
R3608 VGND.n112 VGND.n111 760.639
R3609 VGND.n106 VGND.n105 760.639
R3610 VGND.n100 VGND.n99 760.639
R3611 VGND.n94 VGND.n93 760.639
R3612 VGND.n88 VGND.n85 760.639
R3613 VGND.n1050 VGND.n712 744.222
R3614 VGND.n1025 VGND.n711 744.222
R3615 VGND.n1022 VGND.n713 744.222
R3616 VGND.n334 VGND.n333 744.222
R3617 VGND.n1738 VGND.n337 744.222
R3618 VGND.n1042 VGND.n1033 744.222
R3619 VGND.n1128 VGND.n581 744.222
R3620 VGND.n589 VGND.n580 744.222
R3621 VGND.n586 VGND.n583 744.222
R3622 VGND.n1115 VGND.n603 744.222
R3623 VGND.n613 VGND.n602 744.222
R3624 VGND.n610 VGND.n604 744.222
R3625 VGND.n1102 VGND.n627 744.222
R3626 VGND.n637 VGND.n626 744.222
R3627 VGND.n634 VGND.n628 744.222
R3628 VGND.n1089 VGND.n651 744.222
R3629 VGND.n661 VGND.n650 744.222
R3630 VGND.n658 VGND.n652 744.222
R3631 VGND.n1076 VGND.n675 744.222
R3632 VGND.n685 VGND.n674 744.222
R3633 VGND.n682 VGND.n676 744.222
R3634 VGND.n717 VGND.n716 744.222
R3635 VGND.n718 VGND.n699 744.222
R3636 VGND.n1071 VGND.n695 744.222
R3637 VGND.n1252 VGND.n1251 742.855
R3638 VGND.n1231 VGND.n1230 742.855
R3639 VGND.n1367 VGND.n1366 742.855
R3640 VGND.n1342 VGND.n1341 742.855
R3641 VGND.n1317 VGND.n1316 742.855
R3642 VGND.n1292 VGND.n1291 742.855
R3643 VGND.n1204 VGND.n1203 742.855
R3644 VGND.n1185 VGND.n553 742.855
R3645 VGND.n1252 VGND.n552 719.461
R3646 VGND.n1231 VGND.n551 719.461
R3647 VGND.n1367 VGND.n550 719.461
R3648 VGND.n1342 VGND.n549 719.461
R3649 VGND.n1317 VGND.n548 719.461
R3650 VGND.n1292 VGND.n547 719.461
R3651 VGND.n1203 VGND.n546 719.461
R3652 VGND.n1718 VGND.n553 719.461
R3653 VGND.n1601 VGND.n1599 631.795
R3654 VGND.n1692 VGND.n1691 631.795
R3655 VGND.n1625 VGND.n1623 631.795
R3656 VGND.n1674 VGND.n1673 631.795
R3657 VGND.n1652 VGND.n1650 631.795
R3658 VGND.n1656 VGND.n1655 631.795
R3659 VGND.n728 VGND.t562 607.409
R3660 VGND.n171 VGND.t563 607.409
R3661 VGND.n1035 VGND.n1032 587.761
R3662 VGND.n1744 VGND.n1743 587.761
R3663 VGND.n1021 VGND.n714 587.761
R3664 VGND.n1027 VGND.n710 587.761
R3665 VGND.n681 VGND.n677 587.761
R3666 VGND.n687 VGND.n673 587.761
R3667 VGND.n657 VGND.n653 587.761
R3668 VGND.n663 VGND.n649 587.761
R3669 VGND.n633 VGND.n629 587.761
R3670 VGND.n639 VGND.n625 587.761
R3671 VGND.n609 VGND.n605 587.761
R3672 VGND.n615 VGND.n601 587.761
R3673 VGND.n585 VGND.n584 587.761
R3674 VGND.n591 VGND.n579 587.761
R3675 VGND.n697 VGND.n694 587.761
R3676 VGND.n724 VGND.n723 587.761
R3677 VGND.n725 VGND.n724 585
R3678 VGND.n698 VGND.n697 585
R3679 VGND.n688 VGND.n687 585
R3680 VGND.n681 VGND.n680 585
R3681 VGND.n664 VGND.n663 585
R3682 VGND.n657 VGND.n656 585
R3683 VGND.n640 VGND.n639 585
R3684 VGND.n633 VGND.n632 585
R3685 VGND.n616 VGND.n615 585
R3686 VGND.n609 VGND.n608 585
R3687 VGND.n592 VGND.n591 585
R3688 VGND.n585 VGND.n564 585
R3689 VGND.n1745 VGND.n1744 585
R3690 VGND.n1036 VGND.n1035 585
R3691 VGND.n1028 VGND.n1027 585
R3692 VGND.n1021 VGND.n1020 585
R3693 VGND.n1235 VGND.n538 561.451
R3694 VGND.n1385 VGND.n539 561.451
R3695 VGND.n1375 VGND.n540 561.451
R3696 VGND.n1350 VGND.n541 561.451
R3697 VGND.n1325 VGND.n542 561.451
R3698 VGND.n1300 VGND.n543 561.451
R3699 VGND.n1176 VGND.n544 561.451
R3700 VGND.n1720 VGND.n536 561.451
R3701 VGND.n1597 VGND.t521 549.061
R3702 VGND.t13 VGND.n1597 549.061
R3703 VGND.n1599 VGND.t6 549.061
R3704 VGND.t121 VGND.n1601 549.061
R3705 VGND.n1602 VGND.t493 549.061
R3706 VGND.t268 VGND.n1602 549.061
R3707 VGND.n1692 VGND.t266 549.061
R3708 VGND.n1691 VGND.t506 549.061
R3709 VGND.n1621 VGND.t502 549.061
R3710 VGND.t280 VGND.n1621 549.061
R3711 VGND.n1623 VGND.t495 549.061
R3712 VGND.t115 VGND.n1625 549.061
R3713 VGND.n1626 VGND.t188 549.061
R3714 VGND.t299 VGND.n1626 549.061
R3715 VGND.n1674 VGND.t428 549.061
R3716 VGND.n1673 VGND.t117 549.061
R3717 VGND.n1648 VGND.t278 549.061
R3718 VGND.t252 VGND.n1648 549.061
R3719 VGND.n1650 VGND.t213 549.061
R3720 VGND.t558 VGND.n1652 549.061
R3721 VGND.n1653 VGND.t430 549.061
R3722 VGND.t421 VGND.n1653 549.061
R3723 VGND.n1656 VGND.t423 549.061
R3724 VGND.n1655 VGND.t380 549.061
R3725 VGND.n1795 VGND.t371 549.061
R3726 VGND.n1795 VGND.t363 549.061
R3727 VGND.n1187 VGND.n552 541.75
R3728 VGND.n1219 VGND.n551 541.75
R3729 VGND.n1190 VGND.n550 541.75
R3730 VGND.n1216 VGND.n549 541.75
R3731 VGND.n1193 VGND.n548 541.75
R3732 VGND.n1213 VGND.n547 541.75
R3733 VGND.n1196 VGND.n546 541.75
R3734 VGND.n1718 VGND.n535 541.75
R3735 VGND.n1023 VGND.n1022 540.784
R3736 VGND.n1023 VGND.n711 540.784
R3737 VGND.n1039 VGND.n1033 540.784
R3738 VGND.n1039 VGND.n337 540.784
R3739 VGND.n587 VGND.n586 540.784
R3740 VGND.n587 VGND.n580 540.784
R3741 VGND.n611 VGND.n610 540.784
R3742 VGND.n611 VGND.n602 540.784
R3743 VGND.n635 VGND.n634 540.784
R3744 VGND.n635 VGND.n626 540.784
R3745 VGND.n659 VGND.n658 540.784
R3746 VGND.n659 VGND.n650 540.784
R3747 VGND.n683 VGND.n682 540.784
R3748 VGND.n683 VGND.n674 540.784
R3749 VGND.n1068 VGND.n695 540.784
R3750 VGND.n1068 VGND.n699 540.784
R3751 VGND.n1053 VGND.n711 534.99
R3752 VGND.n1053 VGND.n712 534.99
R3753 VGND.n1741 VGND.n337 534.99
R3754 VGND.n1741 VGND.n333 534.99
R3755 VGND.n1131 VGND.n580 534.99
R3756 VGND.n1131 VGND.n581 534.99
R3757 VGND.n1118 VGND.n602 534.99
R3758 VGND.n1118 VGND.n603 534.99
R3759 VGND.n1105 VGND.n626 534.99
R3760 VGND.n1105 VGND.n627 534.99
R3761 VGND.n1092 VGND.n650 534.99
R3762 VGND.n1092 VGND.n651 534.99
R3763 VGND.n1079 VGND.n674 534.99
R3764 VGND.n1079 VGND.n675 534.99
R3765 VGND.n721 VGND.n699 534.99
R3766 VGND.n721 VGND.n717 534.99
R3767 VGND.n1187 VGND.n538 507.276
R3768 VGND.n1219 VGND.n539 507.276
R3769 VGND.n1190 VGND.n540 507.276
R3770 VGND.n1216 VGND.n541 507.276
R3771 VGND.n1193 VGND.n542 507.276
R3772 VGND.n1213 VGND.n543 507.276
R3773 VGND.n1196 VGND.n544 507.276
R3774 VGND.n1720 VGND.n535 507.276
R3775 VGND.t489 VGND.t146 491.372
R3776 VGND.t294 VGND.t489 491.372
R3777 VGND.t457 VGND.t294 491.372
R3778 VGND.t290 VGND.t417 491.372
R3779 VGND.t288 VGND.t290 491.372
R3780 VGND.t419 VGND.t288 491.372
R3781 VGND.t150 VGND.t333 491.372
R3782 VGND.t166 VGND.t150 491.372
R3783 VGND.t498 VGND.t166 491.372
R3784 VGND.t207 VGND.t209 491.372
R3785 VGND.t529 VGND.t207 491.372
R3786 VGND.t75 VGND.t529 491.372
R3787 VGND.t350 VGND.t196 491.372
R3788 VGND.t196 VGND.t246 491.372
R3789 VGND.t246 VGND.t352 491.372
R3790 VGND.t340 VGND.t361 491.372
R3791 VGND.t361 VGND.t43 491.372
R3792 VGND.t43 VGND.t338 491.372
R3793 VGND.t519 VGND.t134 491.372
R3794 VGND.t134 VGND.t356 491.372
R3795 VGND.t356 VGND.t136 491.372
R3796 VGND.t69 VGND.t326 491.372
R3797 VGND.t326 VGND.t106 491.372
R3798 VGND.t106 VGND.t104 491.372
R3799 VGND.t447 VGND.t276 491.372
R3800 VGND.t276 VGND.t248 491.372
R3801 VGND.t248 VGND.t152 491.372
R3802 VGND.t388 VGND.t382 491.372
R3803 VGND.t382 VGND.t384 491.372
R3804 VGND.t384 VGND.t386 491.372
R3805 VGND.t408 VGND.t410 491.372
R3806 VGND.t410 VGND.t412 491.372
R3807 VGND.t412 VGND.t414 491.372
R3808 VGND.t272 VGND.t314 491.372
R3809 VGND.t314 VGND.t297 491.372
R3810 VGND.t297 VGND.t312 491.372
R3811 VGND.t310 VGND.t354 491.372
R3812 VGND.t354 VGND.t54 491.372
R3813 VGND.t54 VGND.t52 491.372
R3814 VGND.t17 VGND.t15 491.372
R3815 VGND.t15 VGND.t10 491.372
R3816 VGND.t10 VGND.t19 491.372
R3817 VGND.t556 VGND.t455 491.372
R3818 VGND.t455 VGND.t466 491.372
R3819 VGND.t466 VGND.t119 491.372
R3820 VGND.t440 VGND.t464 491.372
R3821 VGND.t464 VGND.t318 491.372
R3822 VGND.t318 VGND.t211 491.372
R3823 VGND.t100 VGND.t65 491.372
R3824 VGND.t435 VGND.t100 491.372
R3825 VGND.t79 VGND.t435 491.372
R3826 VGND.t102 VGND.t67 471.786
R3827 VGND.n314 VGND.n136 455.522
R3828 VGND.n1003 VGND.n159 442.918
R3829 VGND.n263 VGND.n189 430.216
R3830 VGND.n259 VGND.t0 377.098
R3831 VGND.n227 VGND.t0 377.098
R3832 VGND.n1253 VGND.n1252 356.277
R3833 VGND.n1232 VGND.n1231 356.277
R3834 VGND.n1368 VGND.n1367 356.277
R3835 VGND.n1343 VGND.n1342 356.277
R3836 VGND.n1318 VGND.n1317 356.277
R3837 VGND.n1293 VGND.n1292 356.277
R3838 VGND.n1203 VGND.n1202 356.277
R3839 VGND.n1714 VGND.n553 356.277
R3840 VGND.t56 VGND.n555 346.868
R3841 VGND.n1708 VGND.t127 346.868
R3842 VGND.n261 VGND.n255 334.05
R3843 VGND.t521 VGND.t139 330.94
R3844 VGND.t516 VGND.t13 330.94
R3845 VGND.t527 VGND.t516 330.94
R3846 VGND.t6 VGND.t527 330.94
R3847 VGND.t274 VGND.t121 330.94
R3848 VGND.t533 VGND.t274 330.94
R3849 VGND.t493 VGND.t533 330.94
R3850 VGND.t453 VGND.t268 330.94
R3851 VGND.t270 VGND.t453 330.94
R3852 VGND.t266 VGND.t270 330.94
R3853 VGND.t227 VGND.t506 330.94
R3854 VGND.t504 VGND.t227 330.94
R3855 VGND.t502 VGND.t504 330.94
R3856 VGND.t322 VGND.t280 330.94
R3857 VGND.t123 VGND.t322 330.94
R3858 VGND.t495 VGND.t123 330.94
R3859 VGND.t198 VGND.t115 330.94
R3860 VGND.t330 VGND.t198 330.94
R3861 VGND.t188 VGND.t330 330.94
R3862 VGND.t445 VGND.t299 330.94
R3863 VGND.t443 VGND.t445 330.94
R3864 VGND.t428 VGND.t443 330.94
R3865 VGND.t308 VGND.t117 330.94
R3866 VGND.t491 VGND.t308 330.94
R3867 VGND.t278 VGND.t491 330.94
R3868 VGND.t77 VGND.t252 330.94
R3869 VGND.t552 VGND.t77 330.94
R3870 VGND.t213 VGND.t552 330.94
R3871 VGND.t47 VGND.t558 330.94
R3872 VGND.t523 VGND.t47 330.94
R3873 VGND.t430 VGND.t523 330.94
R3874 VGND.t176 VGND.t421 330.94
R3875 VGND.t174 VGND.t176 330.94
R3876 VGND.t423 VGND.t174 330.94
R3877 VGND.t380 VGND.t374 330.94
R3878 VGND.t374 VGND.t377 330.94
R3879 VGND.t377 VGND.t371 330.94
R3880 VGND.t363 VGND.t365 330.94
R3881 VGND.t8 VGND.n138 325.082
R3882 VGND.t8 VGND.n1760 325.082
R3883 VGND.n728 VGND.t344 321.423
R3884 VGND.n171 VGND.t342 321.423
R3885 VGND.n1791 VGND.n80 303.616
R3886 VGND.n510 VGND.n344 297.553
R3887 VGND.n345 VGND.n344 297.553
R3888 VGND.n363 VGND.n345 297.553
R3889 VGND.n508 VGND.n363 297.553
R3890 VGND.n508 VGND.n364 297.553
R3891 VGND.n364 VGND.n346 297.553
R3892 VGND.n381 VGND.n346 297.553
R3893 VGND.n381 VGND.n362 297.553
R3894 VGND.n387 VGND.n362 297.553
R3895 VGND.n387 VGND.n347 297.553
R3896 VGND.n393 VGND.n347 297.553
R3897 VGND.n393 VGND.n361 297.553
R3898 VGND.n399 VGND.n361 297.553
R3899 VGND.n399 VGND.n348 297.553
R3900 VGND.n405 VGND.n348 297.553
R3901 VGND.n405 VGND.n360 297.553
R3902 VGND.n411 VGND.n360 297.553
R3903 VGND.n411 VGND.n349 297.553
R3904 VGND.n417 VGND.n349 297.553
R3905 VGND.n417 VGND.n359 297.553
R3906 VGND.n423 VGND.n359 297.553
R3907 VGND.n423 VGND.n350 297.553
R3908 VGND.n429 VGND.n350 297.553
R3909 VGND.n429 VGND.n358 297.553
R3910 VGND.n435 VGND.n358 297.553
R3911 VGND.n435 VGND.n351 297.553
R3912 VGND.n441 VGND.n351 297.553
R3913 VGND.n441 VGND.n357 297.553
R3914 VGND.n447 VGND.n357 297.553
R3915 VGND.n447 VGND.n352 297.553
R3916 VGND.n453 VGND.n352 297.553
R3917 VGND.n453 VGND.n356 297.553
R3918 VGND.n459 VGND.n356 297.553
R3919 VGND.n459 VGND.n353 297.553
R3920 VGND.n465 VGND.n353 297.553
R3921 VGND.n465 VGND.n355 297.553
R3922 VGND.n355 VGND.n16 297.553
R3923 VGND.n1823 VGND.n16 297.553
R3924 VGND.n1823 VGND.n17 297.553
R3925 VGND.n17 VGND.n7 297.553
R3926 VGND.n25 VGND.n7 297.553
R3927 VGND.n25 VGND.n15 297.553
R3928 VGND.n31 VGND.n15 297.553
R3929 VGND.n31 VGND.n8 297.553
R3930 VGND.n37 VGND.n8 297.553
R3931 VGND.n37 VGND.n14 297.553
R3932 VGND.n43 VGND.n14 297.553
R3933 VGND.n43 VGND.n9 297.553
R3934 VGND.n49 VGND.n9 297.553
R3935 VGND.n49 VGND.n13 297.553
R3936 VGND.n55 VGND.n13 297.553
R3937 VGND.n55 VGND.n10 297.553
R3938 VGND.n61 VGND.n10 297.553
R3939 VGND.n61 VGND.n12 297.553
R3940 VGND.n1790 VGND.n85 297.553
R3941 VGND.n85 VGND.n76 297.553
R3942 VGND.n93 VGND.n76 297.553
R3943 VGND.n93 VGND.n83 297.553
R3944 VGND.n99 VGND.n83 297.553
R3945 VGND.n99 VGND.n77 297.553
R3946 VGND.n105 VGND.n77 297.553
R3947 VGND.n105 VGND.n82 297.553
R3948 VGND.n111 VGND.n82 297.553
R3949 VGND.n111 VGND.n78 297.553
R3950 VGND.n117 VGND.n78 297.553
R3951 VGND.n117 VGND.n81 297.553
R3952 VGND.n123 VGND.n81 297.553
R3953 VGND.n123 VGND.n79 297.553
R3954 VGND.n158 VGND.n142 292.5
R3955 VGND.n771 VGND.n158 292.5
R3956 VGND.n1751 VGND.n162 292.5
R3957 VGND.n771 VGND.n162 292.5
R3958 VGND.n228 VGND.n225 292.5
R3959 VGND.n262 VGND.n225 292.5
R3960 VGND.n223 VGND.n222 292.5
R3961 VGND.n262 VGND.n223 292.5
R3962 VGND.n858 VGND.n165 288.961
R3963 VGND.n1759 VGND.n141 288.961
R3964 VGND.n258 VGND.n216 288.961
R3965 VGND.n252 VGND.n251 288.961
R3966 VGND.n263 VGND.t346 285.123
R3967 VGND.n1236 VGND.n1235 281.135
R3968 VGND.n1386 VGND.n1385 281.135
R3969 VGND.n1376 VGND.n1375 281.135
R3970 VGND.n1351 VGND.n1350 281.135
R3971 VGND.n1326 VGND.n1325 281.135
R3972 VGND.n1301 VGND.n1300 281.135
R3973 VGND.n1176 VGND.n519 281.135
R3974 VGND.n536 VGND.n529 281.135
R3975 VGND.t365 VGND.t367 275.329
R3976 VGND.n262 VGND.n261 258.13
R3977 VGND.n1001 VGND.n999 257.264
R3978 VGND.n151 VGND.t132 254.272
R3979 VGND.t139 VGND.t200 246.464
R3980 VGND.n565 VGND.t163 230.401
R3981 VGND.n1036 VGND.n1034 226.917
R3982 VGND.n1750 VGND.n165 223.68
R3983 VGND.n1759 VGND.n1758 223.68
R3984 VGND.n258 VGND.n257 223.68
R3985 VGND.n253 VGND.n252 223.68
R3986 VGND.n1763 VGND.n1762 220.702
R3987 VGND.t67 VGND.t302 209.071
R3988 VGND.t302 VGND.t56 209.071
R3989 VGND.t200 VGND.t127 209.071
R3990 VGND.n858 VGND.n163 205.69
R3991 VGND.n156 VGND.n141 205.69
R3992 VGND.n266 VGND.n216 205.69
R3993 VGND.n251 VGND.n232 205.69
R3994 VGND.n1728 VGND.n514 200.744
R3995 VGND.n1303 VGND.n1302 200.744
R3996 VGND.n1328 VGND.n1327 200.744
R3997 VGND.n1353 VGND.n1352 200.744
R3998 VGND.n1378 VGND.n1377 200.744
R3999 VGND.n1387 VGND.n1223 200.744
R4000 VGND.n1260 VGND.n1237 200.744
R4001 VGND.n1724 VGND.n1723 200.744
R4002 VGND.n1028 VGND.n166 196.581
R4003 VGND.n1793 VGND.n1792 195.292
R4004 VGND.n89 VGND.n88 195
R4005 VGND.n88 VGND.n80 195
R4006 VGND.n95 VGND.n94 195
R4007 VGND.n94 VGND.n80 195
R4008 VGND.n101 VGND.n100 195
R4009 VGND.n100 VGND.n80 195
R4010 VGND.n107 VGND.n106 195
R4011 VGND.n106 VGND.n80 195
R4012 VGND.n113 VGND.n112 195
R4013 VGND.n112 VGND.n80 195
R4014 VGND.n119 VGND.n118 195
R4015 VGND.n118 VGND.n80 195
R4016 VGND.n125 VGND.n124 195
R4017 VGND.n124 VGND.n80 195
R4018 VGND.n1774 VGND.n1773 195
R4019 VGND.n1773 VGND.n80 195
R4020 VGND.n86 VGND.n84 195
R4021 VGND.n84 VGND.n80 195
R4022 VGND.n21 VGND.n20 195
R4023 VGND.n20 VGND.n11 195
R4024 VGND.n27 VGND.n26 195
R4025 VGND.n26 VGND.n11 195
R4026 VGND.n33 VGND.n32 195
R4027 VGND.n32 VGND.n11 195
R4028 VGND.n39 VGND.n38 195
R4029 VGND.n38 VGND.n11 195
R4030 VGND.n45 VGND.n44 195
R4031 VGND.n44 VGND.n11 195
R4032 VGND.n51 VGND.n50 195
R4033 VGND.n50 VGND.n11 195
R4034 VGND.n57 VGND.n56 195
R4035 VGND.n56 VGND.n11 195
R4036 VGND.n63 VGND.n62 195
R4037 VGND.n62 VGND.n11 195
R4038 VGND.n1805 VGND.n1804 195
R4039 VGND.n1804 VGND.n11 195
R4040 VGND.n369 VGND.n368 195
R4041 VGND.n368 VGND.n354 195
R4042 VGND.n367 VGND.n366 195
R4043 VGND.n366 VGND.n354 195
R4044 VGND.n377 VGND.n376 195
R4045 VGND.n376 VGND.n354 195
R4046 VGND.n383 VGND.n382 195
R4047 VGND.n382 VGND.n354 195
R4048 VGND.n389 VGND.n388 195
R4049 VGND.n388 VGND.n354 195
R4050 VGND.n395 VGND.n394 195
R4051 VGND.n394 VGND.n354 195
R4052 VGND.n401 VGND.n400 195
R4053 VGND.n400 VGND.n354 195
R4054 VGND.n407 VGND.n406 195
R4055 VGND.n406 VGND.n354 195
R4056 VGND.n413 VGND.n412 195
R4057 VGND.n412 VGND.n354 195
R4058 VGND.n419 VGND.n418 195
R4059 VGND.n418 VGND.n354 195
R4060 VGND.n425 VGND.n424 195
R4061 VGND.n424 VGND.n354 195
R4062 VGND.n431 VGND.n430 195
R4063 VGND.n430 VGND.n354 195
R4064 VGND.n437 VGND.n436 195
R4065 VGND.n436 VGND.n354 195
R4066 VGND.n443 VGND.n442 195
R4067 VGND.n442 VGND.n354 195
R4068 VGND.n449 VGND.n448 195
R4069 VGND.n448 VGND.n354 195
R4070 VGND.n455 VGND.n454 195
R4071 VGND.n454 VGND.n354 195
R4072 VGND.n461 VGND.n460 195
R4073 VGND.n460 VGND.n354 195
R4074 VGND.n467 VGND.n466 195
R4075 VGND.n466 VGND.n354 195
R4076 VGND.n471 VGND.n470 195
R4077 VGND.n470 VGND.n354 195
R4078 VGND.n343 VGND.n340 195
R4079 VGND.n354 VGND.n343 195
R4080 VGND.n872 VGND.n752 195
R4081 VGND.n990 VGND.n752 195
R4082 VGND.n854 VGND.n753 195
R4083 VGND.n990 VGND.n753 195
R4084 VGND.n877 VGND.n751 195
R4085 VGND.n990 VGND.n751 195
R4086 VGND.n851 VGND.n754 195
R4087 VGND.n990 VGND.n754 195
R4088 VGND.n894 VGND.n750 195
R4089 VGND.n990 VGND.n750 195
R4090 VGND.n840 VGND.n755 195
R4091 VGND.n990 VGND.n755 195
R4092 VGND.n899 VGND.n749 195
R4093 VGND.n990 VGND.n749 195
R4094 VGND.n837 VGND.n756 195
R4095 VGND.n990 VGND.n756 195
R4096 VGND.n916 VGND.n748 195
R4097 VGND.n990 VGND.n748 195
R4098 VGND.n826 VGND.n757 195
R4099 VGND.n990 VGND.n757 195
R4100 VGND.n921 VGND.n747 195
R4101 VGND.n990 VGND.n747 195
R4102 VGND.n823 VGND.n758 195
R4103 VGND.n990 VGND.n758 195
R4104 VGND.n938 VGND.n746 195
R4105 VGND.n990 VGND.n746 195
R4106 VGND.n812 VGND.n759 195
R4107 VGND.n990 VGND.n759 195
R4108 VGND.n943 VGND.n745 195
R4109 VGND.n990 VGND.n745 195
R4110 VGND.n809 VGND.n760 195
R4111 VGND.n990 VGND.n760 195
R4112 VGND.n960 VGND.n744 195
R4113 VGND.n990 VGND.n744 195
R4114 VGND.n798 VGND.n761 195
R4115 VGND.n990 VGND.n761 195
R4116 VGND.n965 VGND.n743 195
R4117 VGND.n990 VGND.n743 195
R4118 VGND.n795 VGND.n762 195
R4119 VGND.n990 VGND.n762 195
R4120 VGND.n765 VGND.n742 195
R4121 VGND.n990 VGND.n742 195
R4122 VGND.n988 VGND.n987 195
R4123 VGND.n990 VGND.n988 195
R4124 VGND.n992 VGND.n991 195
R4125 VGND.n991 VGND.n990 195
R4126 VGND.n989 VGND.n738 195
R4127 VGND.n990 VGND.n989 195
R4128 VGND.n150 VGND.n149 195
R4129 VGND.n151 VGND.n150 195
R4130 VGND.n153 VGND.n152 195
R4131 VGND.n152 VGND.n151 195
R4132 VGND.n243 VGND.n242 195
R4133 VGND.n242 VGND.n241 195
R4134 VGND.n240 VGND.n235 195
R4135 VGND.n241 VGND.n240 195
R4136 VGND.n272 VGND.n207 195
R4137 VGND.n301 VGND.n207 195
R4138 VGND.n213 VGND.n209 195
R4139 VGND.n301 VGND.n209 195
R4140 VGND.n212 VGND.n206 195
R4141 VGND.n301 VGND.n206 195
R4142 VGND.n281 VGND.n280 195
R4143 VGND.n301 VGND.n281 195
R4144 VGND.n291 VGND.n205 195
R4145 VGND.n301 VGND.n205 195
R4146 VGND.n286 VGND.n282 195
R4147 VGND.n301 VGND.n282 195
R4148 VGND.n285 VGND.n204 195
R4149 VGND.n301 VGND.n204 195
R4150 VGND.n300 VGND.n299 195
R4151 VGND.n301 VGND.n300 195
R4152 VGND.t367 VGND.t369 191.115
R4153 VGND.n186 VGND.n184 190.601
R4154 VGND.n1209 VGND.n1208 184.73
R4155 VGND.n1299 VGND.n1285 184.73
R4156 VGND.n1324 VGND.n1310 184.73
R4157 VGND.n1349 VGND.n1335 184.73
R4158 VGND.n1374 VGND.n1360 184.73
R4159 VGND.n1390 VGND.n1389 184.73
R4160 VGND.n1247 VGND.n1246 184.73
R4161 VGND.n1722 VGND.n533 184.73
R4162 VGND VGND.n728 161.595
R4163 VGND VGND.n171 161.595
R4164 VGND.n1726 VGND.n524 155.677
R4165 VGND.n1728 VGND.n517 152.744
R4166 VGND.n1303 VGND.n1277 152.744
R4167 VGND.n1328 VGND.n1274 152.744
R4168 VGND.n1353 VGND.n1271 152.744
R4169 VGND.n1378 VGND.n1268 152.744
R4170 VGND.n1234 VGND.n1223 152.744
R4171 VGND.n1260 VGND.n1259 152.744
R4172 VGND.n1724 VGND.n530 152.744
R4173 VGND.t369 VGND.n1794 149.852
R4174 VGND.n509 VGND.n354 146.72
R4175 VGND.n1534 VGND.n1523 146.25
R4176 VGND.n1535 VGND.n1534 146.25
R4177 VGND.n1545 VGND.n1544 146.25
R4178 VGND.n1546 VGND.n1545 146.25
R4179 VGND.n1411 VGND.n1410 146.25
R4180 VGND.n1410 VGND.n1409 146.25
R4181 VGND.n1419 VGND.n1412 146.25
R4182 VGND.n1420 VGND.n1419 146.25
R4183 VGND.n1511 VGND.n1423 146.25
R4184 VGND.n1423 VGND.n1422 146.25
R4185 VGND.n1431 VGND.n1424 146.25
R4186 VGND.n1432 VGND.n1431 146.25
R4187 VGND.n1502 VGND.n1435 146.25
R4188 VGND.n1435 VGND.n1434 146.25
R4189 VGND.n1443 VGND.n1436 146.25
R4190 VGND.n1444 VGND.n1443 146.25
R4191 VGND.n1493 VGND.n1447 146.25
R4192 VGND.n1447 VGND.n1446 146.25
R4193 VGND.n1455 VGND.n1448 146.25
R4194 VGND.n1456 VGND.n1455 146.25
R4195 VGND.n1484 VGND.n1459 146.25
R4196 VGND.n1459 VGND.n1458 146.25
R4197 VGND.n1467 VGND.n1460 146.25
R4198 VGND.n1468 VGND.n1467 146.25
R4199 VGND.n1475 VGND.n1471 146.25
R4200 VGND.n1471 VGND.n1470 146.25
R4201 VGND.n1552 VGND.n1551 146.25
R4202 VGND.n1551 VGND.n1550 146.25
R4203 VGND.n1160 VGND.n1150 146.25
R4204 VGND.n1161 VGND.n1160 146.25
R4205 VGND.n1149 VGND.n1148 146.25
R4206 VGND.n1148 VGND.n1147 146.25
R4207 VGND.n1566 VGND.n1565 146.25
R4208 VGND.n1567 VGND.n1566 146.25
R4209 VGND.n1707 VGND.n1706 146.25
R4210 VGND.n1708 VGND.n1707 146.25
R4211 VGND.n1532 VGND.n1531 146.25
R4212 VGND.n1532 VGND.n555 146.25
R4213 VGND.n1654 VGND.n74 146.25
R4214 VGND.n1655 VGND.n1654 146.25
R4215 VGND.n1658 VGND.n1657 146.25
R4216 VGND.n1657 VGND.n1656 146.25
R4217 VGND.n1651 VGND.n1634 146.25
R4218 VGND.n1652 VGND.n1651 146.25
R4219 VGND.n1649 VGND.n1633 146.25
R4220 VGND.n1650 VGND.n1649 146.25
R4221 VGND.n1672 VGND.n1671 146.25
R4222 VGND.n1673 VGND.n1672 146.25
R4223 VGND.n1676 VGND.n1675 146.25
R4224 VGND.n1675 VGND.n1674 146.25
R4225 VGND.n1624 VGND.n1610 146.25
R4226 VGND.n1625 VGND.n1624 146.25
R4227 VGND.n1622 VGND.n1609 146.25
R4228 VGND.n1623 VGND.n1622 146.25
R4229 VGND.n1690 VGND.n1689 146.25
R4230 VGND.n1691 VGND.n1690 146.25
R4231 VGND.n1694 VGND.n1693 146.25
R4232 VGND.n1693 VGND.n1692 146.25
R4233 VGND.n1600 VGND.n1586 146.25
R4234 VGND.n1601 VGND.n1600 146.25
R4235 VGND.n1598 VGND.n1585 146.25
R4236 VGND.n1599 VGND.n1598 146.25
R4237 VGND.n1792 VGND.n69 146.25
R4238 VGND.n1775 VGND.n79 146.25
R4239 VGND.n1791 VGND.n79 146.25
R4240 VGND.n1777 VGND.n81 146.25
R4241 VGND.n1791 VGND.n81 146.25
R4242 VGND.n1779 VGND.n78 146.25
R4243 VGND.n1791 VGND.n78 146.25
R4244 VGND.n1781 VGND.n82 146.25
R4245 VGND.n1791 VGND.n82 146.25
R4246 VGND.n1783 VGND.n77 146.25
R4247 VGND.n1791 VGND.n77 146.25
R4248 VGND.n1785 VGND.n83 146.25
R4249 VGND.n1791 VGND.n83 146.25
R4250 VGND.n1787 VGND.n76 146.25
R4251 VGND.n1791 VGND.n76 146.25
R4252 VGND.n1790 VGND.n1789 146.25
R4253 VGND.n1791 VGND.n1790 146.25
R4254 VGND.n1806 VGND.n12 146.25
R4255 VGND.n1824 VGND.n12 146.25
R4256 VGND.n1808 VGND.n10 146.25
R4257 VGND.n1824 VGND.n10 146.25
R4258 VGND.n1810 VGND.n13 146.25
R4259 VGND.n1824 VGND.n13 146.25
R4260 VGND.n1812 VGND.n9 146.25
R4261 VGND.n1824 VGND.n9 146.25
R4262 VGND.n1814 VGND.n14 146.25
R4263 VGND.n1824 VGND.n14 146.25
R4264 VGND.n1816 VGND.n8 146.25
R4265 VGND.n1824 VGND.n8 146.25
R4266 VGND.n1818 VGND.n15 146.25
R4267 VGND.n1824 VGND.n15 146.25
R4268 VGND.n1820 VGND.n7 146.25
R4269 VGND.n1824 VGND.n7 146.25
R4270 VGND.n1823 VGND.n1822 146.25
R4271 VGND.n1824 VGND.n1823 146.25
R4272 VGND.n475 VGND.n355 146.25
R4273 VGND.n509 VGND.n355 146.25
R4274 VGND.n477 VGND.n353 146.25
R4275 VGND.n509 VGND.n353 146.25
R4276 VGND.n479 VGND.n356 146.25
R4277 VGND.n509 VGND.n356 146.25
R4278 VGND.n481 VGND.n352 146.25
R4279 VGND.n509 VGND.n352 146.25
R4280 VGND.n483 VGND.n357 146.25
R4281 VGND.n509 VGND.n357 146.25
R4282 VGND.n485 VGND.n351 146.25
R4283 VGND.n509 VGND.n351 146.25
R4284 VGND.n487 VGND.n358 146.25
R4285 VGND.n509 VGND.n358 146.25
R4286 VGND.n489 VGND.n350 146.25
R4287 VGND.n509 VGND.n350 146.25
R4288 VGND.n491 VGND.n359 146.25
R4289 VGND.n509 VGND.n359 146.25
R4290 VGND.n493 VGND.n349 146.25
R4291 VGND.n509 VGND.n349 146.25
R4292 VGND.n495 VGND.n360 146.25
R4293 VGND.n509 VGND.n360 146.25
R4294 VGND.n497 VGND.n348 146.25
R4295 VGND.n509 VGND.n348 146.25
R4296 VGND.n499 VGND.n361 146.25
R4297 VGND.n509 VGND.n361 146.25
R4298 VGND.n501 VGND.n347 146.25
R4299 VGND.n509 VGND.n347 146.25
R4300 VGND.n503 VGND.n362 146.25
R4301 VGND.n509 VGND.n362 146.25
R4302 VGND.n505 VGND.n346 146.25
R4303 VGND.n509 VGND.n346 146.25
R4304 VGND.n508 VGND.n507 146.25
R4305 VGND.n509 VGND.n508 146.25
R4306 VGND.n371 VGND.n345 146.25
R4307 VGND.n509 VGND.n345 146.25
R4308 VGND.n511 VGND.n510 146.25
R4309 VGND.n510 VGND.n509 146.25
R4310 VGND.n1756 VGND.n1755 146.25
R4311 VGND.n1755 VGND.n1754 146.25
R4312 VGND.n1753 VGND.n1752 146.25
R4313 VGND.n1754 VGND.n1753 146.25
R4314 VGND.n873 VGND.n856 146.25
R4315 VGND.n856 VGND.n771 146.25
R4316 VGND.n878 VGND.n853 146.25
R4317 VGND.n853 VGND.n771 146.25
R4318 VGND.n882 VGND.n780 146.25
R4319 VGND.n976 VGND.n780 146.25
R4320 VGND.n846 VGND.n782 146.25
R4321 VGND.n976 VGND.n782 146.25
R4322 VGND.n888 VGND.n779 146.25
R4323 VGND.n976 VGND.n779 146.25
R4324 VGND.n843 VGND.n783 146.25
R4325 VGND.n976 VGND.n783 146.25
R4326 VGND.n895 VGND.n842 146.25
R4327 VGND.n842 VGND.n771 146.25
R4328 VGND.n900 VGND.n839 146.25
R4329 VGND.n839 VGND.n771 146.25
R4330 VGND.n904 VGND.n778 146.25
R4331 VGND.n976 VGND.n778 146.25
R4332 VGND.n832 VGND.n784 146.25
R4333 VGND.n976 VGND.n784 146.25
R4334 VGND.n910 VGND.n777 146.25
R4335 VGND.n976 VGND.n777 146.25
R4336 VGND.n829 VGND.n785 146.25
R4337 VGND.n976 VGND.n785 146.25
R4338 VGND.n917 VGND.n828 146.25
R4339 VGND.n828 VGND.n771 146.25
R4340 VGND.n922 VGND.n825 146.25
R4341 VGND.n825 VGND.n771 146.25
R4342 VGND.n926 VGND.n776 146.25
R4343 VGND.n976 VGND.n776 146.25
R4344 VGND.n818 VGND.n786 146.25
R4345 VGND.n976 VGND.n786 146.25
R4346 VGND.n932 VGND.n775 146.25
R4347 VGND.n976 VGND.n775 146.25
R4348 VGND.n815 VGND.n787 146.25
R4349 VGND.n976 VGND.n787 146.25
R4350 VGND.n939 VGND.n814 146.25
R4351 VGND.n814 VGND.n771 146.25
R4352 VGND.n944 VGND.n811 146.25
R4353 VGND.n811 VGND.n771 146.25
R4354 VGND.n948 VGND.n774 146.25
R4355 VGND.n976 VGND.n774 146.25
R4356 VGND.n804 VGND.n788 146.25
R4357 VGND.n976 VGND.n788 146.25
R4358 VGND.n954 VGND.n773 146.25
R4359 VGND.n976 VGND.n773 146.25
R4360 VGND.n801 VGND.n789 146.25
R4361 VGND.n976 VGND.n789 146.25
R4362 VGND.n961 VGND.n800 146.25
R4363 VGND.n800 VGND.n771 146.25
R4364 VGND.n966 VGND.n797 146.25
R4365 VGND.n797 VGND.n771 146.25
R4366 VGND.n794 VGND.n772 146.25
R4367 VGND.n976 VGND.n772 146.25
R4368 VGND.n974 VGND.n973 146.25
R4369 VGND.n976 VGND.n974 146.25
R4370 VGND.n978 VGND.n977 146.25
R4371 VGND.n977 VGND.n976 146.25
R4372 VGND.n975 VGND.n766 146.25
R4373 VGND.n976 VGND.n975 146.25
R4374 VGND.n764 VGND.n763 146.25
R4375 VGND.n771 VGND.n763 146.25
R4376 VGND.n993 VGND.n740 146.25
R4377 VGND.n771 VGND.n740 146.25
R4378 VGND.n1007 VGND.n1006 146.25
R4379 VGND.n1006 VGND.n1005 146.25
R4380 VGND.n1000 VGND.n733 146.25
R4381 VGND.n1001 VGND.n1000 146.25
R4382 VGND.n998 VGND.n732 146.25
R4383 VGND.n999 VGND.n998 146.25
R4384 VGND.n1016 VGND.n1015 146.25
R4385 VGND.n1017 VGND.n1016 146.25
R4386 VGND.n145 VGND.n144 146.25
R4387 VGND.n146 VGND.n145 146.25
R4388 VGND.n244 VGND.n237 146.25
R4389 VGND.n238 VGND.n237 146.25
R4390 VGND.n231 VGND.n224 146.25
R4391 VGND.n263 VGND.n224 146.25
R4392 VGND.n265 VGND.n264 146.25
R4393 VGND.n264 VGND.n263 146.25
R4394 VGND.n273 VGND.n215 146.25
R4395 VGND.n215 VGND.n191 146.25
R4396 VGND.n211 VGND.n210 146.25
R4397 VGND.n210 VGND.n191 146.25
R4398 VGND.n305 VGND.n304 146.25
R4399 VGND.n304 VGND.n303 146.25
R4400 VGND.n302 VGND.n199 146.25
R4401 VGND.n303 VGND.n302 146.25
R4402 VGND.n195 VGND.n193 146.25
R4403 VGND.n303 VGND.n193 146.25
R4404 VGND.n194 VGND.n192 146.25
R4405 VGND.n303 VGND.n192 146.25
R4406 VGND.n292 VGND.n288 146.25
R4407 VGND.n288 VGND.n191 146.25
R4408 VGND.n284 VGND.n283 146.25
R4409 VGND.n283 VGND.n191 146.25
R4410 VGND.n319 VGND.n318 146.25
R4411 VGND.n318 VGND.n317 146.25
R4412 VGND.n185 VGND.n176 146.25
R4413 VGND.n186 VGND.n185 146.25
R4414 VGND.n183 VGND.n175 146.25
R4415 VGND.n184 VGND.n183 146.25
R4416 VGND.n328 VGND.n327 146.25
R4417 VGND.n329 VGND.n328 146.25
R4418 VGND.n1751 VGND.n1750 143.361
R4419 VGND.n1758 VGND.n142 143.361
R4420 VGND.n257 VGND.n222 143.361
R4421 VGND.n253 VGND.n228 143.361
R4422 VGND.n606 VGND.n592 141.846
R4423 VGND.n630 VGND.n616 141.846
R4424 VGND.n654 VGND.n640 141.846
R4425 VGND.n678 VGND.n664 141.846
R4426 VGND.n696 VGND.n688 141.846
R4427 VGND.n315 VGND.n314 141.596
R4428 VGND.n608 VGND.n606 141.343
R4429 VGND.n632 VGND.n630 141.343
R4430 VGND.n656 VGND.n654 141.343
R4431 VGND.n680 VGND.n678 141.343
R4432 VGND.n698 VGND.n696 141.343
R4433 VGND.n1005 VGND.n1004 140.327
R4434 VGND.t304 VGND.n208 135.933
R4435 VGND.n1020 VGND.n1018 135.099
R4436 VGND.n1797 VGND.n69 133.755
R4437 VGND.n1797 VGND.n74 133.755
R4438 VGND.n1659 VGND.n1658 133.755
R4439 VGND.n1659 VGND.n1634 133.755
R4440 VGND.n1633 VGND.n1628 133.755
R4441 VGND.n1671 VGND.n1628 133.755
R4442 VGND.n1677 VGND.n1676 133.755
R4443 VGND.n1677 VGND.n1610 133.755
R4444 VGND.n1609 VGND.n1604 133.755
R4445 VGND.n1689 VGND.n1604 133.755
R4446 VGND.n1695 VGND.n1694 133.755
R4447 VGND.n1695 VGND.n1586 133.755
R4448 VGND.n1585 VGND.n1580 133.755
R4449 VGND.n1706 VGND.n1580 133.755
R4450 VGND.n1538 VGND.n1531 133.755
R4451 VGND.n1538 VGND.n1523 133.755
R4452 VGND.n1544 VGND.n1402 133.755
R4453 VGND.n1411 VGND.n1402 133.755
R4454 VGND.n1512 VGND.n1412 133.755
R4455 VGND.n1512 VGND.n1511 133.755
R4456 VGND.n1503 VGND.n1424 133.755
R4457 VGND.n1503 VGND.n1502 133.755
R4458 VGND.n1494 VGND.n1436 133.755
R4459 VGND.n1494 VGND.n1493 133.755
R4460 VGND.n1485 VGND.n1448 133.755
R4461 VGND.n1485 VGND.n1484 133.755
R4462 VGND.n1476 VGND.n1460 133.755
R4463 VGND.n1476 VGND.n1475 133.755
R4464 VGND.n1553 VGND.n1552 133.755
R4465 VGND.n1553 VGND.n1150 133.755
R4466 VGND.n1149 VGND.n567 133.755
R4467 VGND.n1565 VGND.n567 133.755
R4468 VGND.n241 VGND.n239 133.377
R4469 VGND.n1211 VGND.n1210 131.84
R4470 VGND.n1287 VGND.n1286 131.84
R4471 VGND.n1312 VGND.n1311 131.84
R4472 VGND.n1337 VGND.n1336 131.84
R4473 VGND.n1362 VGND.n1361 131.84
R4474 VGND.n1392 VGND.n1391 131.84
R4475 VGND.n1248 VGND.n1242 131.84
R4476 VGND.n1397 VGND.n1396 131.84
R4477 VGND.n1206 VGND.n1205 125.35
R4478 VGND.n1289 VGND.n1288 125.35
R4479 VGND.n1314 VGND.n1313 125.35
R4480 VGND.n1339 VGND.n1338 125.35
R4481 VGND.n1364 VGND.n1363 125.35
R4482 VGND.n1229 VGND.n1222 125.35
R4483 VGND.n1250 VGND.n1249 125.35
R4484 VGND.n1398 VGND.n554 125.35
R4485 VGND.n255 VGND.t0 123.16
R4486 VGND.n313 VGND.n191 118.132
R4487 VGND.n1715 VGND.n1714 117.001
R4488 VGND.n1714 VGND.n1713 117.001
R4489 VGND.n1202 VGND.n1201 117.001
R4490 VGND.n1202 VGND.n545 117.001
R4491 VGND.n1207 VGND.n544 117.001
R4492 VGND.n1719 VGND.n544 117.001
R4493 VGND.n1294 VGND.n1293 117.001
R4494 VGND.n1293 VGND.n545 117.001
R4495 VGND.n1298 VGND.n543 117.001
R4496 VGND.n1719 VGND.n543 117.001
R4497 VGND.n1319 VGND.n1318 117.001
R4498 VGND.n1318 VGND.n545 117.001
R4499 VGND.n1323 VGND.n542 117.001
R4500 VGND.n1719 VGND.n542 117.001
R4501 VGND.n1344 VGND.n1343 117.001
R4502 VGND.n1343 VGND.n545 117.001
R4503 VGND.n1348 VGND.n541 117.001
R4504 VGND.n1719 VGND.n541 117.001
R4505 VGND.n1369 VGND.n1368 117.001
R4506 VGND.n1368 VGND.n545 117.001
R4507 VGND.n1373 VGND.n540 117.001
R4508 VGND.n1719 VGND.n540 117.001
R4509 VGND.n1233 VGND.n1232 117.001
R4510 VGND.n1232 VGND.n545 117.001
R4511 VGND.n1388 VGND.n539 117.001
R4512 VGND.n1719 VGND.n539 117.001
R4513 VGND.n1254 VGND.n1253 117.001
R4514 VGND.n1253 VGND.n545 117.001
R4515 VGND.n1245 VGND.n538 117.001
R4516 VGND.n1719 VGND.n538 117.001
R4517 VGND.n1721 VGND.n1720 117.001
R4518 VGND.n1720 VGND.n1719 117.001
R4519 VGND.t426 VGND.t98 115.859
R4520 VGND.n1824 VGND.n11 114.246
R4521 VGND.n1017 VGND.t459 112.261
R4522 VGND.n999 VGND.t345 112.261
R4523 VGND.t90 VGND.n1001 112.261
R4524 VGND.n1005 VGND.t396 112.261
R4525 VGND.n1211 VGND.n1198 111.68
R4526 VGND.n1297 VGND.n1286 111.68
R4527 VGND.n1322 VGND.n1311 111.68
R4528 VGND.n1347 VGND.n1336 111.68
R4529 VGND.n1372 VGND.n1361 111.68
R4530 VGND.n1392 VGND.n1221 111.68
R4531 VGND.n1244 VGND.n1242 111.68
R4532 VGND.n1396 VGND.n534 111.68
R4533 VGND.n1710 VGND.n1709 111.663
R4534 VGND.n1833 VGND.n1 110.933
R4535 VGND.n1833 VGND.n1832 110.933
R4536 VGND.n1765 VGND.n130 110.933
R4537 VGND.n1765 VGND.n132 110.933
R4538 VGND.n320 VGND.n176 105.695
R4539 VGND.n320 VGND.n319 105.695
R4540 VGND.n311 VGND.n194 105.695
R4541 VGND.n311 VGND.n195 105.695
R4542 VGND.n306 VGND.n199 105.695
R4543 VGND.n306 VGND.n305 105.695
R4544 VGND.n1008 VGND.n733 105.695
R4545 VGND.n1008 VGND.n1007 105.695
R4546 VGND.n979 VGND.n766 105.695
R4547 VGND.n979 VGND.n978 105.695
R4548 VGND.n973 VGND.n791 105.695
R4549 VGND.n794 VGND.n791 105.695
R4550 VGND.n955 VGND.n801 105.695
R4551 VGND.n955 VGND.n954 105.695
R4552 VGND.n949 VGND.n804 105.695
R4553 VGND.n949 VGND.n948 105.695
R4554 VGND.n933 VGND.n815 105.695
R4555 VGND.n933 VGND.n932 105.695
R4556 VGND.n927 VGND.n818 105.695
R4557 VGND.n927 VGND.n926 105.695
R4558 VGND.n911 VGND.n829 105.695
R4559 VGND.n911 VGND.n910 105.695
R4560 VGND.n905 VGND.n832 105.695
R4561 VGND.n905 VGND.n904 105.695
R4562 VGND.n889 VGND.n843 105.695
R4563 VGND.n889 VGND.n888 105.695
R4564 VGND.n883 VGND.n846 105.695
R4565 VGND.n883 VGND.n882 105.695
R4566 VGND.n732 VGND.n727 105.695
R4567 VGND.n1015 VGND.n727 105.695
R4568 VGND.n175 VGND.n170 105.695
R4569 VGND.n327 VGND.n170 105.695
R4570 VGND.n317 VGND.n316 103.965
R4571 VGND.n1794 VGND.t141 102.638
R4572 VGND.n1201 VGND.n517 101.555
R4573 VGND.n1294 VGND.n1277 101.555
R4574 VGND.n1319 VGND.n1274 101.555
R4575 VGND.n1344 VGND.n1271 101.555
R4576 VGND.n1369 VGND.n1268 101.555
R4577 VGND.n1234 VGND.n1233 101.555
R4578 VGND.n1259 VGND.n1254 101.555
R4579 VGND.n1715 VGND.n530 101.555
R4580 VGND.n1004 VGND.n1003 99.0083
R4581 VGND.n1199 VGND.n546 97.5005
R4582 VGND.n1719 VGND.n546 97.5005
R4583 VGND.n1206 VGND.n1178 97.5005
R4584 VGND.n1400 VGND.n1178 97.5005
R4585 VGND.n1209 VGND.n1177 97.5005
R4586 VGND.n1400 VGND.n1177 97.5005
R4587 VGND.n1296 VGND.n547 97.5005
R4588 VGND.n1719 VGND.n547 97.5005
R4589 VGND.n1288 VGND.n1179 97.5005
R4590 VGND.n1400 VGND.n1179 97.5005
R4591 VGND.n1285 VGND.n1175 97.5005
R4592 VGND.n1400 VGND.n1175 97.5005
R4593 VGND.n1321 VGND.n548 97.5005
R4594 VGND.n1719 VGND.n548 97.5005
R4595 VGND.n1313 VGND.n1180 97.5005
R4596 VGND.n1400 VGND.n1180 97.5005
R4597 VGND.n1310 VGND.n1174 97.5005
R4598 VGND.n1400 VGND.n1174 97.5005
R4599 VGND.n1346 VGND.n549 97.5005
R4600 VGND.n1719 VGND.n549 97.5005
R4601 VGND.n1338 VGND.n1181 97.5005
R4602 VGND.n1400 VGND.n1181 97.5005
R4603 VGND.n1335 VGND.n1173 97.5005
R4604 VGND.n1400 VGND.n1173 97.5005
R4605 VGND.n1371 VGND.n550 97.5005
R4606 VGND.n1719 VGND.n550 97.5005
R4607 VGND.n1363 VGND.n1182 97.5005
R4608 VGND.n1400 VGND.n1182 97.5005
R4609 VGND.n1360 VGND.n1172 97.5005
R4610 VGND.n1400 VGND.n1172 97.5005
R4611 VGND.n1227 VGND.n551 97.5005
R4612 VGND.n1719 VGND.n551 97.5005
R4613 VGND.n1222 VGND.n1183 97.5005
R4614 VGND.n1400 VGND.n1183 97.5005
R4615 VGND.n1390 VGND.n1171 97.5005
R4616 VGND.n1400 VGND.n1171 97.5005
R4617 VGND.n1243 VGND.n552 97.5005
R4618 VGND.n1719 VGND.n552 97.5005
R4619 VGND.n1249 VGND.n1184 97.5005
R4620 VGND.n1400 VGND.n1184 97.5005
R4621 VGND.n1247 VGND.n1170 97.5005
R4622 VGND.n1400 VGND.n1170 97.5005
R4623 VGND.n1718 VGND.n1717 97.5005
R4624 VGND.n1719 VGND.n1718 97.5005
R4625 VGND.n1399 VGND.n1398 97.5005
R4626 VGND.n1400 VGND.n1399 97.5005
R4627 VGND.n1169 VGND.n533 97.5005
R4628 VGND.n1400 VGND.n1169 97.5005
R4629 VGND.n134 VGND.n130 97.5005
R4630 VGND.n1762 VGND.n134 97.5005
R4631 VGND.n133 VGND.n132 97.5005
R4632 VGND.n1762 VGND.n133 97.5005
R4633 VGND.n1832 VGND.n1831 97.5005
R4634 VGND.n1831 VGND.n1830 97.5005
R4635 VGND.n1829 VGND.n1 97.5005
R4636 VGND.n1830 VGND.n1829 97.5005
R4637 VGND.n1752 VGND.n1751 93.4405
R4638 VGND.n1756 VGND.n142 93.4405
R4639 VGND.n265 VGND.n222 93.4405
R4640 VGND.n231 VGND.n228 93.4405
R4641 VGND.n1794 VGND.n1793 93.0698
R4642 VGND.n1400 VGND.n1168 90.9633
R4643 VGND.n1825 VGND.n6 87.9761
R4644 VGND.n1735 VGND.t549 84.5161
R4645 VGND.n1045 VGND.t110 84.5161
R4646 VGND.n1030 VGND.t477 84.5161
R4647 VGND.n1058 VGND.t257 84.5161
R4648 VGND.n1063 VGND.t112 84.5161
R4649 VGND.n701 VGND.t283 84.5161
R4650 VGND.n690 VGND.t216 84.5161
R4651 VGND.n1084 VGND.t192 84.5161
R4652 VGND.n666 VGND.t510 84.5161
R4653 VGND.n1097 VGND.t532 84.5161
R4654 VGND.n642 VGND.t325 84.5161
R4655 VGND.n1110 VGND.t126 84.5161
R4656 VGND.n618 VGND.t555 84.5161
R4657 VGND.n1123 VGND.t321 84.5161
R4658 VGND.n594 VGND.t64 84.5161
R4659 VGND.n1136 VGND.t241 84.5161
R4660 VGND.n236 VGND.t547 84.1574
R4661 VGND.n214 VGND.t399 84.1574
R4662 VGND.n277 VGND.t512 84.1574
R4663 VGND.n287 VGND.t406 84.1574
R4664 VGND.n296 VGND.t305 84.1574
R4665 VGND.n147 VGND.t133 84.1574
R4666 VGND.n855 VGND.t439 84.1574
R4667 VGND.n852 VGND.t258 84.1574
R4668 VGND.n841 VGND.t482 84.1574
R4669 VGND.n838 VGND.t475 84.1574
R4670 VGND.n827 VGND.t264 84.1574
R4671 VGND.n824 VGND.t265 84.1574
R4672 VGND.n813 VGND.t154 84.1574
R4673 VGND.n810 VGND.t89 84.1574
R4674 VGND.n799 VGND.t526 84.1574
R4675 VGND.n796 VGND.t138 84.1574
R4676 VGND.n984 VGND.t407 84.1574
R4677 VGND.n739 VGND.t307 84.1574
R4678 VGND.n129 VGND.t511 84.1574
R4679 VGND.n126 VGND.t262 84.1574
R4680 VGND.n120 VGND.t260 84.1574
R4681 VGND.n114 VGND.t263 84.1574
R4682 VGND.n108 VGND.t261 84.1574
R4683 VGND.n102 VGND.t373 84.1574
R4684 VGND.n96 VGND.t379 84.1574
R4685 VGND.n90 VGND.t376 84.1574
R4686 VGND.n67 VGND.t544 84.1574
R4687 VGND.n64 VGND.t515 84.1574
R4688 VGND.n58 VGND.t187 84.1574
R4689 VGND.n52 VGND.t142 84.1574
R4690 VGND.n46 VGND.t255 84.1574
R4691 VGND.n40 VGND.t203 84.1574
R4692 VGND.n34 VGND.t348 84.1574
R4693 VGND.n28 VGND.t178 84.1574
R4694 VGND.n22 VGND.t538 84.1574
R4695 VGND.n473 VGND.t540 84.1574
R4696 VGND.n468 VGND.t539 84.1574
R4697 VGND.n462 VGND.t537 84.1574
R4698 VGND.n456 VGND.t37 84.1574
R4699 VGND.n450 VGND.t29 84.1574
R4700 VGND.n444 VGND.t41 84.1574
R4701 VGND.n438 VGND.t32 84.1574
R4702 VGND.n432 VGND.t39 84.1574
R4703 VGND.n426 VGND.t38 84.1574
R4704 VGND.n420 VGND.t40 84.1574
R4705 VGND.n414 VGND.t35 84.1574
R4706 VGND.n408 VGND.t30 84.1574
R4707 VGND.n402 VGND.t250 84.1574
R4708 VGND.n396 VGND.t33 84.1574
R4709 VGND.n390 VGND.t34 84.1574
R4710 VGND.n384 VGND.t97 84.1574
R4711 VGND.n378 VGND.t36 84.1574
R4712 VGND.n373 VGND.t31 84.1574
R4713 VGND.n341 VGND.t42 84.1574
R4714 VGND.n201 VGND.t390 83.7172
R4715 VGND.n197 VGND.t316 83.7172
R4716 VGND.n178 VGND.t392 83.7172
R4717 VGND.n174 VGND.t61 83.7172
R4718 VGND.n848 VGND.t130 83.7172
R4719 VGND.n845 VGND.t535 83.7172
R4720 VGND.n834 VGND.t296 83.7172
R4721 VGND.n831 VGND.t4 83.7172
R4722 VGND.n820 VGND.t62 83.7172
R4723 VGND.n817 VGND.t226 83.7172
R4724 VGND.n806 VGND.t242 83.7172
R4725 VGND.n803 VGND.t223 83.7172
R4726 VGND.n793 VGND.t525 83.7172
R4727 VGND.n768 VGND.t359 83.7172
R4728 VGND.n735 VGND.t397 83.7172
R4729 VGND.n731 VGND.t460 83.7172
R4730 VGND.n716 VGND.n704 83.5719
R4731 VGND.n716 VGND.n715 83.5719
R4732 VGND.n718 VGND.n702 83.5719
R4733 VGND.n719 VGND.n718 83.5719
R4734 VGND.n1072 VGND.n1071 83.5719
R4735 VGND.n1071 VGND.n1070 83.5719
R4736 VGND.n1076 VGND.n1075 83.5719
R4737 VGND.n1077 VGND.n1076 83.5719
R4738 VGND.n685 VGND.n672 83.5719
R4739 VGND.n686 VGND.n685 83.5719
R4740 VGND.n676 VGND.n668 83.5719
R4741 VGND.n679 VGND.n676 83.5719
R4742 VGND.n1089 VGND.n1088 83.5719
R4743 VGND.n1090 VGND.n1089 83.5719
R4744 VGND.n661 VGND.n648 83.5719
R4745 VGND.n662 VGND.n661 83.5719
R4746 VGND.n652 VGND.n644 83.5719
R4747 VGND.n655 VGND.n652 83.5719
R4748 VGND.n1102 VGND.n1101 83.5719
R4749 VGND.n1103 VGND.n1102 83.5719
R4750 VGND.n637 VGND.n624 83.5719
R4751 VGND.n638 VGND.n637 83.5719
R4752 VGND.n628 VGND.n620 83.5719
R4753 VGND.n631 VGND.n628 83.5719
R4754 VGND.n1115 VGND.n1114 83.5719
R4755 VGND.n1116 VGND.n1115 83.5719
R4756 VGND.n613 VGND.n600 83.5719
R4757 VGND.n614 VGND.n613 83.5719
R4758 VGND.n604 VGND.n596 83.5719
R4759 VGND.n607 VGND.n604 83.5719
R4760 VGND.n1128 VGND.n1127 83.5719
R4761 VGND.n1129 VGND.n1128 83.5719
R4762 VGND.n589 VGND.n578 83.5719
R4763 VGND.n590 VGND.n589 83.5719
R4764 VGND.n583 VGND.n574 83.5719
R4765 VGND.n583 VGND.n582 83.5719
R4766 VGND.n335 VGND.n334 83.5719
R4767 VGND.n334 VGND.n332 83.5719
R4768 VGND.n1738 VGND.n1737 83.5719
R4769 VGND.n1739 VGND.n1738 83.5719
R4770 VGND.n1043 VGND.n1042 83.5719
R4771 VGND.n1042 VGND.n1041 83.5719
R4772 VGND.n1050 VGND.n1049 83.5719
R4773 VGND.n1051 VGND.n1050 83.5719
R4774 VGND.n1025 VGND.n709 83.5719
R4775 VGND.n1026 VGND.n1025 83.5719
R4776 VGND.n713 VGND.n705 83.5719
R4777 VGND.n1019 VGND.n713 83.5719
R4778 VGND.n184 VGND.t343 83.1719
R4779 VGND.t545 VGND.n186 83.1719
R4780 VGND.n317 VGND.t391 83.1719
R4781 VGND.n1210 VGND.n1206 78.6829
R4782 VGND.n1288 VGND.n1287 78.6829
R4783 VGND.n1313 VGND.n1312 78.6829
R4784 VGND.n1338 VGND.n1337 78.6829
R4785 VGND.n1363 VGND.n1362 78.6829
R4786 VGND.n1391 VGND.n1222 78.6829
R4787 VGND.n1249 VGND.n1248 78.6829
R4788 VGND.n1398 VGND.n1397 78.6829
R4789 VGND.n1018 VGND.n1017 78.6611
R4790 VGND.n1394 VGND.n545 77.9686
R4791 VGND.n1210 VGND.n1209 77.9299
R4792 VGND.n1287 VGND.n1285 77.9299
R4793 VGND.n1312 VGND.n1310 77.9299
R4794 VGND.n1337 VGND.n1335 77.9299
R4795 VGND.n1362 VGND.n1360 77.9299
R4796 VGND.n1391 VGND.n1390 77.9299
R4797 VGND.n1248 VGND.n1247 77.9299
R4798 VGND.n1397 VGND.n533 77.9299
R4799 VGND.n201 VGND.n200 75.905
R4800 VGND.n197 VGND.n196 75.905
R4801 VGND.n178 VGND.n177 75.905
R4802 VGND.n174 VGND.n173 75.905
R4803 VGND.n848 VGND.n847 75.905
R4804 VGND.n845 VGND.n844 75.905
R4805 VGND.n834 VGND.n833 75.905
R4806 VGND.n831 VGND.n830 75.905
R4807 VGND.n820 VGND.n819 75.905
R4808 VGND.n817 VGND.n816 75.905
R4809 VGND.n806 VGND.n805 75.905
R4810 VGND.n803 VGND.n802 75.905
R4811 VGND.n793 VGND.n792 75.905
R4812 VGND.n768 VGND.n767 75.905
R4813 VGND.n735 VGND.n734 75.905
R4814 VGND.n731 VGND.n730 75.905
R4815 VGND.n1018 VGND.n725 74.8287
R4816 VGND.n316 VGND.n315 73.3531
R4817 VGND.n1205 VGND.n1204 73.1255
R4818 VGND.n1204 VGND.n1168 73.1255
R4819 VGND.n1291 VGND.n1289 73.1255
R4820 VGND.n1291 VGND.n1168 73.1255
R4821 VGND.n1316 VGND.n1314 73.1255
R4822 VGND.n1316 VGND.n1168 73.1255
R4823 VGND.n1341 VGND.n1339 73.1255
R4824 VGND.n1341 VGND.n1168 73.1255
R4825 VGND.n1366 VGND.n1364 73.1255
R4826 VGND.n1366 VGND.n1168 73.1255
R4827 VGND.n1230 VGND.n1229 73.1255
R4828 VGND.n1230 VGND.n1168 73.1255
R4829 VGND.n1251 VGND.n1250 73.1255
R4830 VGND.n1251 VGND.n1168 73.1255
R4831 VGND.n1185 VGND.n554 73.1255
R4832 VGND.n1185 VGND.n1168 73.1255
R4833 VGND.n883 VGND.n850 73.1255
R4834 VGND.n850 VGND.n160 73.1255
R4835 VGND.n889 VGND.n887 73.1255
R4836 VGND.n887 VGND.n160 73.1255
R4837 VGND.n905 VGND.n836 73.1255
R4838 VGND.n836 VGND.n160 73.1255
R4839 VGND.n911 VGND.n909 73.1255
R4840 VGND.n909 VGND.n160 73.1255
R4841 VGND.n927 VGND.n822 73.1255
R4842 VGND.n822 VGND.n160 73.1255
R4843 VGND.n933 VGND.n931 73.1255
R4844 VGND.n931 VGND.n160 73.1255
R4845 VGND.n949 VGND.n808 73.1255
R4846 VGND.n808 VGND.n160 73.1255
R4847 VGND.n955 VGND.n953 73.1255
R4848 VGND.n953 VGND.n160 73.1255
R4849 VGND.n791 VGND.n790 73.1255
R4850 VGND.n790 VGND.n160 73.1255
R4851 VGND.n979 VGND.n770 73.1255
R4852 VGND.n770 VGND.n160 73.1255
R4853 VGND.n1008 VGND.n737 73.1255
R4854 VGND.n1002 VGND.n737 73.1255
R4855 VGND.n727 VGND.n726 73.1255
R4856 VGND.n997 VGND.n726 73.1255
R4857 VGND.n306 VGND.n190 73.1255
R4858 VGND.n313 VGND.n190 73.1255
R4859 VGND.n312 VGND.n311 73.1255
R4860 VGND.n313 VGND.n312 73.1255
R4861 VGND.n320 VGND.n180 73.1255
R4862 VGND.n187 VGND.n180 73.1255
R4863 VGND.n170 VGND.n169 73.1255
R4864 VGND.n182 VGND.n169 73.1255
R4865 VGND.n1712 VGND.t12 71.4713
R4866 VGND.n1752 VGND.n163 69.2272
R4867 VGND.n1756 VGND.n156 69.2272
R4868 VGND.n266 VGND.n265 69.2272
R4869 VGND.n232 VGND.n231 69.2272
R4870 VGND.n303 VGND.n191 68.7758
R4871 VGND.n299 VGND.n284 68.7561
R4872 VGND.n285 VGND.n284 68.7561
R4873 VGND.n292 VGND.n286 68.7561
R4874 VGND.n292 VGND.n291 68.7561
R4875 VGND.n280 VGND.n211 68.7561
R4876 VGND.n212 VGND.n211 68.7561
R4877 VGND.n273 VGND.n213 68.7561
R4878 VGND.n273 VGND.n272 68.7561
R4879 VGND.n244 VGND.n235 68.7561
R4880 VGND.n244 VGND.n243 68.7561
R4881 VGND.n993 VGND.n738 68.7561
R4882 VGND.n993 VGND.n992 68.7561
R4883 VGND.n987 VGND.n764 68.7561
R4884 VGND.n765 VGND.n764 68.7561
R4885 VGND.n966 VGND.n795 68.7561
R4886 VGND.n966 VGND.n965 68.7561
R4887 VGND.n961 VGND.n798 68.7561
R4888 VGND.n961 VGND.n960 68.7561
R4889 VGND.n944 VGND.n809 68.7561
R4890 VGND.n944 VGND.n943 68.7561
R4891 VGND.n939 VGND.n812 68.7561
R4892 VGND.n939 VGND.n938 68.7561
R4893 VGND.n922 VGND.n823 68.7561
R4894 VGND.n922 VGND.n921 68.7561
R4895 VGND.n917 VGND.n826 68.7561
R4896 VGND.n917 VGND.n916 68.7561
R4897 VGND.n900 VGND.n837 68.7561
R4898 VGND.n900 VGND.n899 68.7561
R4899 VGND.n895 VGND.n840 68.7561
R4900 VGND.n895 VGND.n894 68.7561
R4901 VGND.n878 VGND.n851 68.7561
R4902 VGND.n878 VGND.n877 68.7561
R4903 VGND.n873 VGND.n854 68.7561
R4904 VGND.n873 VGND.n872 68.7561
R4905 VGND.n1775 VGND.n1774 68.7561
R4906 VGND.n1789 VGND.n86 68.7561
R4907 VGND.n1806 VGND.n1805 68.7561
R4908 VGND.n511 VGND.n340 68.7561
R4909 VGND.n153 VGND.n144 68.7561
R4910 VGND.n149 VGND.n144 68.7561
R4911 VGND.t221 VGND.t459 68.6043
R4912 VGND.t345 VGND.t461 68.6043
R4913 VGND.t404 VGND.t90 68.6043
R4914 VGND.t396 VGND.t393 68.6043
R4915 VGND.n234 VGND.n233 67.5509
R4916 VGND.n218 VGND.n217 67.5509
R4917 VGND.n862 VGND.n861 67.5509
R4918 VGND.n860 VGND.n859 67.5509
R4919 VGND.n1734 VGND.n339 67.1161
R4920 VGND.n1046 VGND.n1044 67.1161
R4921 VGND.n1031 VGND.n1029 67.1161
R4922 VGND.n1059 VGND.n706 67.1161
R4923 VGND.n1062 VGND.n703 67.1161
R4924 VGND.n693 VGND.n692 67.1161
R4925 VGND.n691 VGND.n689 67.1161
R4926 VGND.n1085 VGND.n669 67.1161
R4927 VGND.n667 VGND.n665 67.1161
R4928 VGND.n1098 VGND.n645 67.1161
R4929 VGND.n643 VGND.n641 67.1161
R4930 VGND.n1111 VGND.n621 67.1161
R4931 VGND.n619 VGND.n617 67.1161
R4932 VGND.n1124 VGND.n597 67.1161
R4933 VGND.n595 VGND.n593 67.1161
R4934 VGND.n1137 VGND.n575 67.1161
R4935 VGND.n1800 VGND.n70 66.9639
R4936 VGND.n1799 VGND.n71 66.9639
R4937 VGND.n73 VGND.n72 66.9639
R4938 VGND.n1643 VGND.n1642 66.9639
R4939 VGND.n1641 VGND.n1640 66.9639
R4940 VGND.n1638 VGND.n1637 66.9639
R4941 VGND.n1661 VGND.n1636 66.9639
R4942 VGND.n1662 VGND.n1635 66.9639
R4943 VGND.n1665 VGND.n1632 66.9639
R4944 VGND.n1666 VGND.n1631 66.9639
R4945 VGND.n1668 VGND.n1630 66.9639
R4946 VGND.n1669 VGND.n1629 66.9639
R4947 VGND.n1617 VGND.n1616 66.9639
R4948 VGND.n1614 VGND.n1613 66.9639
R4949 VGND.n1679 VGND.n1612 66.9639
R4950 VGND.n1680 VGND.n1611 66.9639
R4951 VGND.n1683 VGND.n1608 66.9639
R4952 VGND.n1684 VGND.n1607 66.9639
R4953 VGND.n1686 VGND.n1606 66.9639
R4954 VGND.n1687 VGND.n1605 66.9639
R4955 VGND.n1593 VGND.n1592 66.9639
R4956 VGND.n1590 VGND.n1589 66.9639
R4957 VGND.n1697 VGND.n1588 66.9639
R4958 VGND.n1698 VGND.n1587 66.9639
R4959 VGND.n1701 VGND.n1584 66.9639
R4960 VGND.n1702 VGND.n1583 66.9639
R4961 VGND.n1704 VGND.n1582 66.9639
R4962 VGND.n1705 VGND.n1581 66.9639
R4963 VGND.n1529 VGND.n1528 66.9639
R4964 VGND.n1527 VGND.n1526 66.9639
R4965 VGND.n1540 VGND.n1525 66.9639
R4966 VGND.n1541 VGND.n1524 66.9639
R4967 VGND.n1522 VGND.n1403 66.9639
R4968 VGND.n1521 VGND.n1404 66.9639
R4969 VGND.n1519 VGND.n1405 66.9639
R4970 VGND.n1518 VGND.n1406 66.9639
R4971 VGND.n1515 VGND.n1413 66.9639
R4972 VGND.n1514 VGND.n1414 66.9639
R4973 VGND.n1416 VGND.n1415 66.9639
R4974 VGND.n1509 VGND.n1508 66.9639
R4975 VGND.n1506 VGND.n1425 66.9639
R4976 VGND.n1505 VGND.n1426 66.9639
R4977 VGND.n1428 VGND.n1427 66.9639
R4978 VGND.n1500 VGND.n1499 66.9639
R4979 VGND.n1497 VGND.n1437 66.9639
R4980 VGND.n1496 VGND.n1438 66.9639
R4981 VGND.n1440 VGND.n1439 66.9639
R4982 VGND.n1491 VGND.n1490 66.9639
R4983 VGND.n1488 VGND.n1449 66.9639
R4984 VGND.n1487 VGND.n1450 66.9639
R4985 VGND.n1452 VGND.n1451 66.9639
R4986 VGND.n1482 VGND.n1481 66.9639
R4987 VGND.n1479 VGND.n1461 66.9639
R4988 VGND.n1478 VGND.n1462 66.9639
R4989 VGND.n1464 VGND.n1463 66.9639
R4990 VGND.n1473 VGND.n1472 66.9639
R4991 VGND.n1157 VGND.n1156 66.9639
R4992 VGND.n1154 VGND.n1153 66.9639
R4993 VGND.n1555 VGND.n1152 66.9639
R4994 VGND.n1556 VGND.n1151 66.9639
R4995 VGND.n1559 VGND.n1144 66.9639
R4996 VGND.n1560 VGND.n1143 66.9639
R4997 VGND.n1562 VGND.n1142 66.9639
R4998 VGND.n1563 VGND.n1141 66.9639
R4999 VGND.n252 VGND.n227 65.0005
R5000 VGND.n259 VGND.n258 65.0005
R5001 VGND.n1760 VGND.n1759 65.0005
R5002 VGND.n165 VGND.n138 65.0005
R5003 VGND.n1758 VGND.n140 65.0005
R5004 VGND.n1748 VGND.n140 65.0005
R5005 VGND.n1750 VGND.n1749 65.0005
R5006 VGND.n1749 VGND.n1748 65.0005
R5007 VGND.n254 VGND.n253 65.0005
R5008 VGND.n255 VGND.n254 65.0005
R5009 VGND.n257 VGND.n256 65.0005
R5010 VGND.n256 VGND.n255 65.0005
R5011 VGND.n1019 VGND.t284 61.0779
R5012 VGND.n1041 VGND.t50 61.0779
R5013 VGND.n1713 VGND.t163 59.2465
R5014 VGND.n1026 VGND.t256 58.651
R5015 VGND.t476 VGND.n1026 58.651
R5016 VGND.t171 VGND.n1051 58.651
R5017 VGND.n1739 VGND.t109 58.651
R5018 VGND.t548 VGND.n1739 58.651
R5019 VGND.t328 VGND.n332 58.651
R5020 VGND.n1765 VGND.n1764 58.5005
R5021 VGND.n1764 VGND.n1763 58.5005
R5022 VGND.n1833 VGND.n3 58.5005
R5023 VGND.n239 VGND.n3 58.5005
R5024 VGND.n1754 VGND.n159 57.2454
R5025 VGND.n1713 VGND.t426 56.6133
R5026 VGND.n303 VGND.t204 55.8298
R5027 VGND.n1830 VGND.t546 55.0911
R5028 VGND.n1003 VGND.n135 53.6536
R5029 VGND.t58 VGND.t60 50.8275
R5030 VGND.t343 VGND.t449 50.8275
R5031 VGND.t400 VGND.t545 50.8275
R5032 VGND.t391 VGND.t402 50.8275
R5033 VGND.t346 VGND.n262 50.614
R5034 VGND.n1548 VGND.n1400 50.16
R5035 VGND.n1776 VGND.n125 49.4227
R5036 VGND.n1778 VGND.n119 49.4227
R5037 VGND.n1780 VGND.n113 49.4227
R5038 VGND.n1782 VGND.n107 49.4227
R5039 VGND.n1784 VGND.n101 49.4227
R5040 VGND.n1786 VGND.n95 49.4227
R5041 VGND.n1788 VGND.n89 49.4227
R5042 VGND.n1807 VGND.n63 49.4227
R5043 VGND.n1809 VGND.n57 49.4227
R5044 VGND.n1811 VGND.n51 49.4227
R5045 VGND.n1813 VGND.n45 49.4227
R5046 VGND.n1815 VGND.n39 49.4227
R5047 VGND.n1817 VGND.n33 49.4227
R5048 VGND.n1819 VGND.n27 49.4227
R5049 VGND.n1821 VGND.n21 49.4227
R5050 VGND.n471 VGND.n18 49.4227
R5051 VGND.n476 VGND.n467 49.4227
R5052 VGND.n478 VGND.n461 49.4227
R5053 VGND.n480 VGND.n455 49.4227
R5054 VGND.n482 VGND.n449 49.4227
R5055 VGND.n484 VGND.n443 49.4227
R5056 VGND.n486 VGND.n437 49.4227
R5057 VGND.n488 VGND.n431 49.4227
R5058 VGND.n490 VGND.n425 49.4227
R5059 VGND.n492 VGND.n419 49.4227
R5060 VGND.n494 VGND.n413 49.4227
R5061 VGND.n496 VGND.n407 49.4227
R5062 VGND.n498 VGND.n401 49.4227
R5063 VGND.n500 VGND.n395 49.4227
R5064 VGND.n502 VGND.n389 49.4227
R5065 VGND.n504 VGND.n383 49.4227
R5066 VGND.n506 VGND.n377 49.4227
R5067 VGND.n367 VGND.n365 49.4227
R5068 VGND.n369 VGND.n342 49.4227
R5069 VGND.n1726 VGND.n520 48.8605
R5070 VGND.t98 VGND.n1712 48.7138
R5071 VGND.n1743 VGND.n335 48.3561
R5072 VGND.n1737 VGND.n336 48.3561
R5073 VGND.n1043 VGND.n1032 48.3561
R5074 VGND.n1049 VGND.n710 48.3561
R5075 VGND.n1055 VGND.n709 48.3561
R5076 VGND.n714 VGND.n705 48.3561
R5077 VGND.n723 VGND.n704 48.3561
R5078 VGND.n702 VGND.n700 48.3561
R5079 VGND.n1075 VGND.n673 48.3561
R5080 VGND.n1081 VGND.n672 48.3561
R5081 VGND.n677 VGND.n668 48.3561
R5082 VGND.n1088 VGND.n649 48.3561
R5083 VGND.n1094 VGND.n648 48.3561
R5084 VGND.n653 VGND.n644 48.3561
R5085 VGND.n1101 VGND.n625 48.3561
R5086 VGND.n1107 VGND.n624 48.3561
R5087 VGND.n629 VGND.n620 48.3561
R5088 VGND.n1114 VGND.n601 48.3561
R5089 VGND.n1120 VGND.n600 48.3561
R5090 VGND.n605 VGND.n596 48.3561
R5091 VGND.n1127 VGND.n579 48.3561
R5092 VGND.n1133 VGND.n578 48.3561
R5093 VGND.n584 VGND.n574 48.3561
R5094 VGND.n1072 VGND.n694 48.3561
R5095 VGND.n1205 VGND.n1200 48.2672
R5096 VGND.n1295 VGND.n1289 48.2672
R5097 VGND.n1320 VGND.n1314 48.2672
R5098 VGND.n1345 VGND.n1339 48.2672
R5099 VGND.n1370 VGND.n1364 48.2672
R5100 VGND.n1229 VGND.n1228 48.2672
R5101 VGND.n1250 VGND.n1241 48.2672
R5102 VGND.n1716 VGND.n554 48.2672
R5103 VGND.n329 VGND.n168 46.7844
R5104 VGND.n1200 VGND.n1199 46.7472
R5105 VGND.n1296 VGND.n1295 46.7472
R5106 VGND.n1321 VGND.n1320 46.7472
R5107 VGND.n1346 VGND.n1345 46.7472
R5108 VGND.n1371 VGND.n1370 46.7472
R5109 VGND.n1228 VGND.n1227 46.7472
R5110 VGND.n1243 VGND.n1241 46.7472
R5111 VGND.n1717 VGND.n1716 46.7472
R5112 VGND.n1212 VGND.n1211 45.0005
R5113 VGND.n1394 VGND.n1212 45.0005
R5114 VGND.n1286 VGND.n1215 45.0005
R5115 VGND.n1394 VGND.n1215 45.0005
R5116 VGND.n1311 VGND.n1195 45.0005
R5117 VGND.n1394 VGND.n1195 45.0005
R5118 VGND.n1336 VGND.n1218 45.0005
R5119 VGND.n1394 VGND.n1218 45.0005
R5120 VGND.n1361 VGND.n1192 45.0005
R5121 VGND.n1394 VGND.n1192 45.0005
R5122 VGND.n1393 VGND.n1392 45.0005
R5123 VGND.n1394 VGND.n1393 45.0005
R5124 VGND.n1242 VGND.n1189 45.0005
R5125 VGND.n1394 VGND.n1189 45.0005
R5126 VGND.n1396 VGND.n1395 45.0005
R5127 VGND.n1395 VGND.n1394 45.0005
R5128 VGND.n1022 VGND.n1021 42.4907
R5129 VGND.n1027 VGND.n712 42.4907
R5130 VGND.n1035 VGND.n1033 42.4907
R5131 VGND.n1744 VGND.n333 42.4907
R5132 VGND.n586 VGND.n585 42.4907
R5133 VGND.n591 VGND.n581 42.4907
R5134 VGND.n610 VGND.n609 42.4907
R5135 VGND.n615 VGND.n603 42.4907
R5136 VGND.n634 VGND.n633 42.4907
R5137 VGND.n639 VGND.n627 42.4907
R5138 VGND.n658 VGND.n657 42.4907
R5139 VGND.n663 VGND.n651 42.4907
R5140 VGND.n682 VGND.n681 42.4907
R5141 VGND.n687 VGND.n675 42.4907
R5142 VGND.n697 VGND.n695 42.4907
R5143 VGND.n724 VGND.n717 42.4907
R5144 VGND.n2 VGND.t237 42.0841
R5145 VGND.n1767 VGND.t235 42.0841
R5146 VGND.n234 VGND.t347 41.3938
R5147 VGND.n218 VGND.t480 41.3938
R5148 VGND.n862 VGND.t481 41.3938
R5149 VGND.n860 VGND.t479 41.3938
R5150 VGND.n530 VGND.n528 39.0005
R5151 VGND.n565 VGND.n528 39.0005
R5152 VGND.n518 VGND.n517 39.0005
R5153 VGND.n524 VGND.n518 39.0005
R5154 VGND.n1290 VGND.n1277 39.0005
R5155 VGND.n1290 VGND.n524 39.0005
R5156 VGND.n1315 VGND.n1274 39.0005
R5157 VGND.n1315 VGND.n524 39.0005
R5158 VGND.n1340 VGND.n1271 39.0005
R5159 VGND.n1340 VGND.n524 39.0005
R5160 VGND.n1365 VGND.n1268 39.0005
R5161 VGND.n1365 VGND.n524 39.0005
R5162 VGND.n1234 VGND.n1226 39.0005
R5163 VGND.n1226 VGND.n524 39.0005
R5164 VGND.n1259 VGND.n1240 39.0005
R5165 VGND.n1240 VGND.n524 39.0005
R5166 VGND.n141 VGND.n139 39.0005
R5167 VGND.n781 VGND.n139 39.0005
R5168 VGND.n858 VGND.n857 39.0005
R5169 VGND.n857 VGND.n781 39.0005
R5170 VGND.n251 VGND.n226 39.0005
R5171 VGND.n261 VGND.n226 39.0005
R5172 VGND.n260 VGND.n216 39.0005
R5173 VGND.n261 VGND.n260 39.0005
R5174 VGND.n582 VGND.t472 38.0445
R5175 VGND.n607 VGND.t23 38.0445
R5176 VGND.n631 VGND.t513 38.0445
R5177 VGND.n655 VGND.t224 38.0445
R5178 VGND.n679 VGND.t487 38.0445
R5179 VGND.n1070 VGND.t483 38.0445
R5180 VGND.t259 VGND.n80 37.3437
R5181 VGND.n722 VGND.n721 36.563
R5182 VGND.n721 VGND.n720 36.563
R5183 VGND.n1068 VGND.n1067 36.563
R5184 VGND.n1069 VGND.n1068 36.563
R5185 VGND.n1080 VGND.n1079 36.563
R5186 VGND.n1079 VGND.n1078 36.563
R5187 VGND.n683 VGND.n671 36.563
R5188 VGND.n684 VGND.n683 36.563
R5189 VGND.n1093 VGND.n1092 36.563
R5190 VGND.n1092 VGND.n1091 36.563
R5191 VGND.n659 VGND.n647 36.563
R5192 VGND.n660 VGND.n659 36.563
R5193 VGND.n1106 VGND.n1105 36.563
R5194 VGND.n1105 VGND.n1104 36.563
R5195 VGND.n635 VGND.n623 36.563
R5196 VGND.n636 VGND.n635 36.563
R5197 VGND.n1119 VGND.n1118 36.563
R5198 VGND.n1118 VGND.n1117 36.563
R5199 VGND.n611 VGND.n599 36.563
R5200 VGND.n612 VGND.n611 36.563
R5201 VGND.n1132 VGND.n1131 36.563
R5202 VGND.n1131 VGND.n1130 36.563
R5203 VGND.n587 VGND.n577 36.563
R5204 VGND.n588 VGND.n587 36.563
R5205 VGND.n1742 VGND.n1741 36.563
R5206 VGND.n1741 VGND.n1740 36.563
R5207 VGND.n1039 VGND.n1038 36.563
R5208 VGND.n1040 VGND.n1039 36.563
R5209 VGND.n1054 VGND.n1053 36.563
R5210 VGND.n1053 VGND.n1052 36.563
R5211 VGND.n1023 VGND.n708 36.563
R5212 VGND.n1024 VGND.n1023 36.563
R5213 VGND.n590 VGND.t240 36.5328
R5214 VGND.t63 VGND.n590 36.5328
R5215 VGND.t560 VGND.n1129 36.5328
R5216 VGND.n614 VGND.t320 36.5328
R5217 VGND.t554 VGND.n614 36.5328
R5218 VGND.t73 VGND.n1116 36.5328
R5219 VGND.n638 VGND.t125 36.5328
R5220 VGND.t324 VGND.n638 36.5328
R5221 VGND.t205 VGND.n1103 36.5328
R5222 VGND.n662 VGND.t531 36.5328
R5223 VGND.t509 VGND.n662 36.5328
R5224 VGND.t243 VGND.n1090 36.5328
R5225 VGND.n686 VGND.t191 36.5328
R5226 VGND.t215 VGND.n686 36.5328
R5227 VGND.t550 VGND.n1077 36.5328
R5228 VGND.n719 VGND.t282 36.5328
R5229 VGND.t111 VGND.n719 36.5328
R5230 VGND.t485 VGND.n715 36.5328
R5231 VGND.n1208 VGND.n1207 36.4805
R5232 VGND.n1299 VGND.n1298 36.4805
R5233 VGND.n1324 VGND.n1323 36.4805
R5234 VGND.n1349 VGND.n1348 36.4805
R5235 VGND.n1374 VGND.n1373 36.4805
R5236 VGND.n1389 VGND.n1388 36.4805
R5237 VGND.n1246 VGND.n1245 36.4805
R5238 VGND.n1722 VGND.n1721 36.4805
R5239 VGND.t60 VGND.n168 36.388
R5240 VGND.n1719 VGND.n537 35.6059
R5241 VGND.t284 VGND.t229 35.5953
R5242 VGND.t256 VGND.t170 35.5953
R5243 VGND.t286 VGND.t476 35.5953
R5244 VGND.t181 VGND.t171 35.5953
R5245 VGND.t50 VGND.t183 35.5953
R5246 VGND.t332 VGND.t109 35.5953
R5247 VGND.t49 VGND.t548 35.5953
R5248 VGND.t25 VGND.t328 35.5953
R5249 VGND.n1199 VGND.n1198 35.2005
R5250 VGND.n1297 VGND.n1296 35.2005
R5251 VGND.n1322 VGND.n1321 35.2005
R5252 VGND.n1347 VGND.n1346 35.2005
R5253 VGND.n1372 VGND.n1371 35.2005
R5254 VGND.n1227 VGND.n1221 35.2005
R5255 VGND.n1244 VGND.n1243 35.2005
R5256 VGND.n1717 VGND.n534 35.2005
R5257 VGND.n1038 VGND.n1032 35.1378
R5258 VGND.n714 VGND.n708 35.1378
R5259 VGND.n677 VGND.n671 35.1378
R5260 VGND.n653 VGND.n647 35.1378
R5261 VGND.n629 VGND.n623 35.1378
R5262 VGND.n605 VGND.n599 35.1378
R5263 VGND.n584 VGND.n577 35.1378
R5264 VGND.n1067 VGND.n694 35.1378
R5265 VGND.n1038 VGND.n1037 34.7613
R5266 VGND.n1742 VGND.n336 34.7613
R5267 VGND.n1743 VGND.n1742 34.7613
R5268 VGND.n1056 VGND.n708 34.7613
R5269 VGND.n1055 VGND.n1054 34.7613
R5270 VGND.n1054 VGND.n710 34.7613
R5271 VGND.n1082 VGND.n671 34.7613
R5272 VGND.n1081 VGND.n1080 34.7613
R5273 VGND.n1080 VGND.n673 34.7613
R5274 VGND.n1095 VGND.n647 34.7613
R5275 VGND.n1094 VGND.n1093 34.7613
R5276 VGND.n1093 VGND.n649 34.7613
R5277 VGND.n1108 VGND.n623 34.7613
R5278 VGND.n1107 VGND.n1106 34.7613
R5279 VGND.n1106 VGND.n625 34.7613
R5280 VGND.n1121 VGND.n599 34.7613
R5281 VGND.n1120 VGND.n1119 34.7613
R5282 VGND.n1119 VGND.n601 34.7613
R5283 VGND.n1134 VGND.n577 34.7613
R5284 VGND.n1133 VGND.n1132 34.7613
R5285 VGND.n1132 VGND.n579 34.7613
R5286 VGND.n1067 VGND.n1066 34.7613
R5287 VGND.n722 VGND.n700 34.7613
R5288 VGND.n723 VGND.n722 34.7613
R5289 VGND.n997 VGND.t221 34.3024
R5290 VGND.t461 VGND.n997 34.3024
R5291 VGND.n1002 VGND.t404 34.3024
R5292 VGND.t393 VGND.n1002 34.3024
R5293 VGND.n1207 VGND.n1198 32.9605
R5294 VGND.n1298 VGND.n1297 32.9605
R5295 VGND.n1323 VGND.n1322 32.9605
R5296 VGND.n1348 VGND.n1347 32.9605
R5297 VGND.n1373 VGND.n1372 32.9605
R5298 VGND.n1388 VGND.n1221 32.9605
R5299 VGND.n1245 VGND.n1244 32.9605
R5300 VGND.n1721 VGND.n534 32.9605
R5301 VGND.n1282 VGND.t156 31.7728
R5302 VGND.n1307 VGND.t468 31.7728
R5303 VGND.n1332 VGND.t220 31.7728
R5304 VGND.n1357 VGND.t442 31.7728
R5305 VGND.n1382 VGND.t169 31.7728
R5306 VGND.n1264 VGND.t469 31.7728
R5307 VGND.n1257 VGND.t158 31.7728
R5308 VGND.n572 VGND.t164 31.7728
R5309 VGND.n1748 VGND.t88 31.6536
R5310 VGND.n1034 VGND.n166 31.1459
R5311 VGND.n330 VGND.n329 30.6122
R5312 VGND.n1407 VGND.n1402 28.8579
R5313 VGND.n1512 VGND.n1417 28.8579
R5314 VGND.n1503 VGND.n1429 28.8579
R5315 VGND.n1494 VGND.n1441 28.8579
R5316 VGND.n1485 VGND.n1453 28.8579
R5317 VGND.n1476 VGND.n1465 28.8579
R5318 VGND.n1553 VGND.n1155 28.8579
R5319 VGND.n1145 VGND.n567 28.8579
R5320 VGND.n1659 VGND.n1639 28.8579
R5321 VGND.n1647 VGND.n1628 28.8579
R5322 VGND.n1677 VGND.n1615 28.8579
R5323 VGND.n1620 VGND.n1604 28.8579
R5324 VGND.n1695 VGND.n1591 28.8579
R5325 VGND.n1596 VGND.n1580 28.8579
R5326 VGND.n1538 VGND.n1537 28.857
R5327 VGND.n1797 VGND.n1796 28.857
R5328 VGND.n1537 VGND.n1536 28.6936
R5329 VGND.n1796 VGND.n1795 28.6936
R5330 VGND.n1597 VGND.n1596 28.6927
R5331 VGND.n1602 VGND.n1591 28.6927
R5332 VGND.n1621 VGND.n1620 28.6927
R5333 VGND.n1626 VGND.n1615 28.6927
R5334 VGND.n1648 VGND.n1647 28.6927
R5335 VGND.n1653 VGND.n1639 28.6927
R5336 VGND.n1146 VGND.n1145 28.6927
R5337 VGND.n1162 VGND.n1155 28.6927
R5338 VGND.n1469 VGND.n1465 28.6927
R5339 VGND.n1457 VGND.n1453 28.6927
R5340 VGND.n1445 VGND.n1441 28.6927
R5341 VGND.n1433 VGND.n1429 28.6927
R5342 VGND.n1421 VGND.n1417 28.6927
R5343 VGND.n1408 VGND.n1407 28.6927
R5344 VGND.n1746 VGND.n1745 28.3145
R5345 VGND.t204 VGND.n301 26.7015
R5346 VGND.t478 VGND.n160 26.0413
R5347 VGND.n516 VGND.n515 25.9728
R5348 VGND.n1281 VGND.n1280 25.9728
R5349 VGND.n1305 VGND.n1279 25.9728
R5350 VGND.n1306 VGND.n1278 25.9728
R5351 VGND.n1330 VGND.n1276 25.9728
R5352 VGND.n1331 VGND.n1275 25.9728
R5353 VGND.n1355 VGND.n1273 25.9728
R5354 VGND.n1356 VGND.n1272 25.9728
R5355 VGND.n1380 VGND.n1270 25.9728
R5356 VGND.n1381 VGND.n1269 25.9728
R5357 VGND.n1266 VGND.n1224 25.9728
R5358 VGND.n1265 VGND.n1225 25.9728
R5359 VGND.n1239 VGND.n1238 25.9728
R5360 VGND.n1256 VGND.n1255 25.9728
R5361 VGND.n570 VGND.n569 25.9728
R5362 VGND.n571 VGND.n568 25.9728
R5363 VGND.n1733 VGND.n335 25.8532
R5364 VGND.n1737 VGND.n1736 25.8532
R5365 VGND.n1047 VGND.n1043 25.8532
R5366 VGND.n1049 VGND.n1048 25.8532
R5367 VGND.n709 VGND.n707 25.8532
R5368 VGND.n1060 VGND.n705 25.8532
R5369 VGND.n1061 VGND.n704 25.8532
R5370 VGND.n1064 VGND.n702 25.8532
R5371 VGND.n1075 VGND.n1074 25.8532
R5372 VGND.n672 VGND.n670 25.8532
R5373 VGND.n1086 VGND.n668 25.8532
R5374 VGND.n1088 VGND.n1087 25.8532
R5375 VGND.n648 VGND.n646 25.8532
R5376 VGND.n1099 VGND.n644 25.8532
R5377 VGND.n1101 VGND.n1100 25.8532
R5378 VGND.n624 VGND.n622 25.8532
R5379 VGND.n1112 VGND.n620 25.8532
R5380 VGND.n1114 VGND.n1113 25.8532
R5381 VGND.n600 VGND.n598 25.8532
R5382 VGND.n1125 VGND.n596 25.8532
R5383 VGND.n1127 VGND.n1126 25.8532
R5384 VGND.n578 VGND.n576 25.8532
R5385 VGND.n1138 VGND.n574 25.8532
R5386 VGND.n1073 VGND.n1072 25.8532
R5387 VGND.n182 VGND.t58 25.414
R5388 VGND.t449 VGND.n182 25.414
R5389 VGND.n187 VGND.t400 25.414
R5390 VGND.t402 VGND.n187 25.414
R5391 VGND.n157 VGND.n156 24.3755
R5392 VGND.n159 VGND.n157 24.3755
R5393 VGND.n163 VGND.n161 24.3755
R5394 VGND.n161 VGND.n159 24.3755
R5395 VGND.n232 VGND.n230 24.3755
R5396 VGND.n230 VGND.n189 24.3755
R5397 VGND.n266 VGND.n220 24.3755
R5398 VGND.n220 VGND.n189 24.3755
R5399 VGND.n1201 VGND.n1200 23.1494
R5400 VGND.n1295 VGND.n1294 23.1494
R5401 VGND.n1320 VGND.n1319 23.1494
R5402 VGND.n1345 VGND.n1344 23.1494
R5403 VGND.n1370 VGND.n1369 23.1494
R5404 VGND.n1233 VGND.n1228 23.1494
R5405 VGND.n1254 VGND.n1241 23.1494
R5406 VGND.n1716 VGND.n1715 23.1494
R5407 VGND.n1719 VGND.n545 23.131
R5408 VGND.n1302 VGND.n1301 22.5005
R5409 VGND.n1301 VGND.n537 22.5005
R5410 VGND.n1327 VGND.n1326 22.5005
R5411 VGND.n1326 VGND.n537 22.5005
R5412 VGND.n1352 VGND.n1351 22.5005
R5413 VGND.n1351 VGND.n537 22.5005
R5414 VGND.n1377 VGND.n1376 22.5005
R5415 VGND.n1376 VGND.n537 22.5005
R5416 VGND.n1387 VGND.n1386 22.5005
R5417 VGND.n1386 VGND.n537 22.5005
R5418 VGND.n1237 VGND.n1236 22.5005
R5419 VGND.n1236 VGND.n537 22.5005
R5420 VGND.n1723 VGND.n529 22.5005
R5421 VGND.n537 VGND.n529 22.5005
R5422 VGND.n519 VGND.n514 22.5005
R5423 VGND.n1711 VGND.n519 22.5005
R5424 VGND.t472 VGND.t542 22.1718
R5425 VGND.t240 VGND.t193 22.1718
R5426 VGND.t474 VGND.t63 22.1718
R5427 VGND.t84 VGND.t560 22.1718
R5428 VGND.t23 VGND.t336 22.1718
R5429 VGND.t320 VGND.t72 22.1718
R5430 VGND.t22 VGND.t554 22.1718
R5431 VGND.t185 VGND.t73 22.1718
R5432 VGND.t513 VGND.t82 22.1718
R5433 VGND.t125 VGND.t306 22.1718
R5434 VGND.t173 VGND.t324 22.1718
R5435 VGND.t144 VGND.t205 22.1718
R5436 VGND.t224 VGND.t433 22.1718
R5437 VGND.t531 VGND.t508 22.1718
R5438 VGND.t239 VGND.t509 22.1718
R5439 VGND.t179 VGND.t243 22.1718
R5440 VGND.t487 VGND.t148 22.1718
R5441 VGND.t191 VGND.t71 22.1718
R5442 VGND.t293 VGND.t215 22.1718
R5443 VGND.t45 VGND.t550 22.1718
R5444 VGND.t483 VGND.t232 22.1718
R5445 VGND.t282 VGND.t238 22.1718
R5446 VGND.t349 VGND.t111 22.1718
R5447 VGND.t113 VGND.t485 22.1718
R5448 VGND.t12 VGND.n524 20.0123
R5449 VGND.n1712 VGND.n1711 19.4911
R5450 VGND.n1789 VGND.n1788 19.3338
R5451 VGND.n1788 VGND.n1787 19.3338
R5452 VGND.n1787 VGND.n1786 19.3338
R5453 VGND.n1786 VGND.n1785 19.3338
R5454 VGND.n1785 VGND.n1784 19.3338
R5455 VGND.n1784 VGND.n1783 19.3338
R5456 VGND.n1783 VGND.n1782 19.3338
R5457 VGND.n1782 VGND.n1781 19.3338
R5458 VGND.n1781 VGND.n1780 19.3338
R5459 VGND.n1780 VGND.n1779 19.3338
R5460 VGND.n1779 VGND.n1778 19.3338
R5461 VGND.n1778 VGND.n1777 19.3338
R5462 VGND.n1777 VGND.n1776 19.3338
R5463 VGND.n1776 VGND.n1775 19.3338
R5464 VGND.n511 VGND.n342 19.3338
R5465 VGND.n371 VGND.n342 19.3338
R5466 VGND.n371 VGND.n365 19.3338
R5467 VGND.n507 VGND.n365 19.3338
R5468 VGND.n507 VGND.n506 19.3338
R5469 VGND.n506 VGND.n505 19.3338
R5470 VGND.n505 VGND.n504 19.3338
R5471 VGND.n504 VGND.n503 19.3338
R5472 VGND.n503 VGND.n502 19.3338
R5473 VGND.n502 VGND.n501 19.3338
R5474 VGND.n501 VGND.n500 19.3338
R5475 VGND.n500 VGND.n499 19.3338
R5476 VGND.n499 VGND.n498 19.3338
R5477 VGND.n498 VGND.n497 19.3338
R5478 VGND.n497 VGND.n496 19.3338
R5479 VGND.n496 VGND.n495 19.3338
R5480 VGND.n495 VGND.n494 19.3338
R5481 VGND.n494 VGND.n493 19.3338
R5482 VGND.n493 VGND.n492 19.3338
R5483 VGND.n492 VGND.n491 19.3338
R5484 VGND.n491 VGND.n490 19.3338
R5485 VGND.n490 VGND.n489 19.3338
R5486 VGND.n489 VGND.n488 19.3338
R5487 VGND.n488 VGND.n487 19.3338
R5488 VGND.n487 VGND.n486 19.3338
R5489 VGND.n486 VGND.n485 19.3338
R5490 VGND.n485 VGND.n484 19.3338
R5491 VGND.n484 VGND.n483 19.3338
R5492 VGND.n483 VGND.n482 19.3338
R5493 VGND.n482 VGND.n481 19.3338
R5494 VGND.n481 VGND.n480 19.3338
R5495 VGND.n480 VGND.n479 19.3338
R5496 VGND.n479 VGND.n478 19.3338
R5497 VGND.n478 VGND.n477 19.3338
R5498 VGND.n477 VGND.n476 19.3338
R5499 VGND.n476 VGND.n475 19.3338
R5500 VGND.n475 VGND.n18 19.3338
R5501 VGND.n1822 VGND.n18 19.3338
R5502 VGND.n1822 VGND.n1821 19.3338
R5503 VGND.n1821 VGND.n1820 19.3338
R5504 VGND.n1820 VGND.n1819 19.3338
R5505 VGND.n1819 VGND.n1818 19.3338
R5506 VGND.n1818 VGND.n1817 19.3338
R5507 VGND.n1817 VGND.n1816 19.3338
R5508 VGND.n1816 VGND.n1815 19.3338
R5509 VGND.n1815 VGND.n1814 19.3338
R5510 VGND.n1814 VGND.n1813 19.3338
R5511 VGND.n1813 VGND.n1812 19.3338
R5512 VGND.n1812 VGND.n1811 19.3338
R5513 VGND.n1811 VGND.n1810 19.3338
R5514 VGND.n1810 VGND.n1809 19.3338
R5515 VGND.n1809 VGND.n1808 19.3338
R5516 VGND.n1808 VGND.n1807 19.3338
R5517 VGND.n1807 VGND.n1806 19.3338
R5518 VGND.n976 VGND.n771 19.0821
R5519 VGND.t170 VGND.n1024 19.0113
R5520 VGND.n1040 VGND.t332 19.0113
R5521 VGND.n301 VGND.t304 18.6103
R5522 VGND.n1208 VGND.n514 18.2672
R5523 VGND.n1302 VGND.n1299 18.2672
R5524 VGND.n1327 VGND.n1324 18.2672
R5525 VGND.n1352 VGND.n1349 18.2672
R5526 VGND.n1377 VGND.n1374 18.2672
R5527 VGND.n1389 VGND.n1387 18.2672
R5528 VGND.n1246 VGND.n1237 18.2672
R5529 VGND.n1723 VGND.n1722 18.2672
R5530 VGND.n354 VGND.t28 18.0461
R5531 VGND.n1052 VGND.t286 17.7979
R5532 VGND.n1052 VGND.t181 17.7979
R5533 VGND.n1740 VGND.t49 17.7979
R5534 VGND.n1740 VGND.t25 17.7979
R5535 VGND.n233 VGND.t360 17.4005
R5536 VGND.n233 VGND.t432 17.4005
R5537 VGND.n217 VGND.t143 17.4005
R5538 VGND.n217 VGND.t1 17.4005
R5539 VGND.n200 VGND.t395 17.4005
R5540 VGND.n200 VGND.t398 17.4005
R5541 VGND.n196 VGND.t497 17.4005
R5542 VGND.n196 VGND.t245 17.4005
R5543 VGND.n177 VGND.t401 17.4005
R5544 VGND.n177 VGND.t403 17.4005
R5545 VGND.n173 VGND.t59 17.4005
R5546 VGND.n173 VGND.t450 17.4005
R5547 VGND.n861 VGND.t9 17.4005
R5548 VGND.n861 VGND.t416 17.4005
R5549 VGND.n859 VGND.t81 17.4005
R5550 VGND.n859 VGND.t27 17.4005
R5551 VGND.n847 VGND.t131 17.4005
R5552 VGND.n847 VGND.t202 17.4005
R5553 VGND.n844 VGND.t292 17.4005
R5554 VGND.n844 VGND.t536 17.4005
R5555 VGND.n833 VGND.t518 17.4005
R5556 VGND.n833 VGND.t231 17.4005
R5557 VGND.n830 VGND.t5 17.4005
R5558 VGND.n830 VGND.t3 17.4005
R5559 VGND.n819 VGND.t438 17.4005
R5560 VGND.n819 VGND.t437 17.4005
R5561 VGND.n816 VGND.t541 17.4005
R5562 VGND.n816 VGND.t287 17.4005
R5563 VGND.n805 VGND.t500 17.4005
R5564 VGND.n805 VGND.t501 17.4005
R5565 VGND.n802 VGND.t87 17.4005
R5566 VGND.n802 VGND.t86 17.4005
R5567 VGND.n792 VGND.t108 17.4005
R5568 VGND.n792 VGND.t463 17.4005
R5569 VGND.n767 VGND.t358 17.4005
R5570 VGND.n767 VGND.t190 17.4005
R5571 VGND.n734 VGND.t405 17.4005
R5572 VGND.n734 VGND.t394 17.4005
R5573 VGND.n730 VGND.t222 17.4005
R5574 VGND.n730 VGND.t462 17.4005
R5575 VGND.n70 VGND.t368 17.4005
R5576 VGND.n70 VGND.t370 17.4005
R5577 VGND.n71 VGND.t364 17.4005
R5578 VGND.n71 VGND.t366 17.4005
R5579 VGND.n72 VGND.t378 17.4005
R5580 VGND.n72 VGND.t372 17.4005
R5581 VGND.n1642 VGND.t381 17.4005
R5582 VGND.n1642 VGND.t375 17.4005
R5583 VGND.n1640 VGND.t175 17.4005
R5584 VGND.n1640 VGND.t424 17.4005
R5585 VGND.n1637 VGND.t422 17.4005
R5586 VGND.n1637 VGND.t177 17.4005
R5587 VGND.n1636 VGND.t524 17.4005
R5588 VGND.n1636 VGND.t431 17.4005
R5589 VGND.n1635 VGND.t559 17.4005
R5590 VGND.n1635 VGND.t48 17.4005
R5591 VGND.n1632 VGND.t553 17.4005
R5592 VGND.n1632 VGND.t214 17.4005
R5593 VGND.n1631 VGND.t253 17.4005
R5594 VGND.n1631 VGND.t78 17.4005
R5595 VGND.n1630 VGND.t492 17.4005
R5596 VGND.n1630 VGND.t279 17.4005
R5597 VGND.n1629 VGND.t118 17.4005
R5598 VGND.n1629 VGND.t309 17.4005
R5599 VGND.n1616 VGND.t444 17.4005
R5600 VGND.n1616 VGND.t429 17.4005
R5601 VGND.n1613 VGND.t300 17.4005
R5602 VGND.n1613 VGND.t446 17.4005
R5603 VGND.n1612 VGND.t331 17.4005
R5604 VGND.n1612 VGND.t189 17.4005
R5605 VGND.n1611 VGND.t116 17.4005
R5606 VGND.n1611 VGND.t199 17.4005
R5607 VGND.n1608 VGND.t124 17.4005
R5608 VGND.n1608 VGND.t496 17.4005
R5609 VGND.n1607 VGND.t281 17.4005
R5610 VGND.n1607 VGND.t323 17.4005
R5611 VGND.n1606 VGND.t505 17.4005
R5612 VGND.n1606 VGND.t503 17.4005
R5613 VGND.n1605 VGND.t507 17.4005
R5614 VGND.n1605 VGND.t228 17.4005
R5615 VGND.n1592 VGND.t271 17.4005
R5616 VGND.n1592 VGND.t267 17.4005
R5617 VGND.n1589 VGND.t269 17.4005
R5618 VGND.n1589 VGND.t454 17.4005
R5619 VGND.n1588 VGND.t534 17.4005
R5620 VGND.n1588 VGND.t494 17.4005
R5621 VGND.n1587 VGND.t122 17.4005
R5622 VGND.n1587 VGND.t275 17.4005
R5623 VGND.n1584 VGND.t528 17.4005
R5624 VGND.n1584 VGND.t7 17.4005
R5625 VGND.n1583 VGND.t14 17.4005
R5626 VGND.n1583 VGND.t517 17.4005
R5627 VGND.n1582 VGND.t140 17.4005
R5628 VGND.n1582 VGND.t522 17.4005
R5629 VGND.n1581 VGND.t128 17.4005
R5630 VGND.n1581 VGND.t201 17.4005
R5631 VGND.n339 VGND.t26 17.4005
R5632 VGND.n339 VGND.t329 17.4005
R5633 VGND.n1044 VGND.t51 17.4005
R5634 VGND.n1044 VGND.t184 17.4005
R5635 VGND.n1029 VGND.t182 17.4005
R5636 VGND.n1029 VGND.t172 17.4005
R5637 VGND.n706 VGND.t285 17.4005
R5638 VGND.n706 VGND.t230 17.4005
R5639 VGND.n703 VGND.t114 17.4005
R5640 VGND.n703 VGND.t486 17.4005
R5641 VGND.n692 VGND.t484 17.4005
R5642 VGND.n692 VGND.t233 17.4005
R5643 VGND.n689 VGND.t46 17.4005
R5644 VGND.n689 VGND.t551 17.4005
R5645 VGND.n669 VGND.t488 17.4005
R5646 VGND.n669 VGND.t149 17.4005
R5647 VGND.n665 VGND.t180 17.4005
R5648 VGND.n665 VGND.t244 17.4005
R5649 VGND.n645 VGND.t225 17.4005
R5650 VGND.n645 VGND.t434 17.4005
R5651 VGND.n641 VGND.t145 17.4005
R5652 VGND.n641 VGND.t206 17.4005
R5653 VGND.n621 VGND.t514 17.4005
R5654 VGND.n621 VGND.t83 17.4005
R5655 VGND.n617 VGND.t186 17.4005
R5656 VGND.n617 VGND.t74 17.4005
R5657 VGND.n597 VGND.t24 17.4005
R5658 VGND.n597 VGND.t337 17.4005
R5659 VGND.n593 VGND.t85 17.4005
R5660 VGND.n593 VGND.t561 17.4005
R5661 VGND.n575 VGND.t473 17.4005
R5662 VGND.n575 VGND.t543 17.4005
R5663 VGND.n1528 VGND.t303 17.4005
R5664 VGND.n1528 VGND.t57 17.4005
R5665 VGND.n1526 VGND.t103 17.4005
R5666 VGND.n1526 VGND.t68 17.4005
R5667 VGND.n1525 VGND.t436 17.4005
R5668 VGND.n1525 VGND.t80 17.4005
R5669 VGND.n1524 VGND.t66 17.4005
R5670 VGND.n1524 VGND.t101 17.4005
R5671 VGND.n1403 VGND.t319 17.4005
R5672 VGND.n1403 VGND.t212 17.4005
R5673 VGND.n1404 VGND.t441 17.4005
R5674 VGND.n1404 VGND.t465 17.4005
R5675 VGND.n1405 VGND.t467 17.4005
R5676 VGND.n1405 VGND.t120 17.4005
R5677 VGND.n1406 VGND.t557 17.4005
R5678 VGND.n1406 VGND.t456 17.4005
R5679 VGND.n1413 VGND.t11 17.4005
R5680 VGND.n1413 VGND.t20 17.4005
R5681 VGND.n1414 VGND.t18 17.4005
R5682 VGND.n1414 VGND.t16 17.4005
R5683 VGND.n1415 VGND.t55 17.4005
R5684 VGND.n1415 VGND.t53 17.4005
R5685 VGND.n1508 VGND.t311 17.4005
R5686 VGND.n1508 VGND.t355 17.4005
R5687 VGND.n1425 VGND.t298 17.4005
R5688 VGND.n1425 VGND.t313 17.4005
R5689 VGND.n1426 VGND.t273 17.4005
R5690 VGND.n1426 VGND.t315 17.4005
R5691 VGND.n1427 VGND.t413 17.4005
R5692 VGND.n1427 VGND.t415 17.4005
R5693 VGND.n1499 VGND.t409 17.4005
R5694 VGND.n1499 VGND.t411 17.4005
R5695 VGND.n1437 VGND.t385 17.4005
R5696 VGND.n1437 VGND.t387 17.4005
R5697 VGND.n1438 VGND.t389 17.4005
R5698 VGND.n1438 VGND.t383 17.4005
R5699 VGND.n1439 VGND.t249 17.4005
R5700 VGND.n1439 VGND.t153 17.4005
R5701 VGND.n1490 VGND.t448 17.4005
R5702 VGND.n1490 VGND.t277 17.4005
R5703 VGND.n1449 VGND.t107 17.4005
R5704 VGND.n1449 VGND.t105 17.4005
R5705 VGND.n1450 VGND.t70 17.4005
R5706 VGND.n1450 VGND.t327 17.4005
R5707 VGND.n1451 VGND.t357 17.4005
R5708 VGND.n1451 VGND.t137 17.4005
R5709 VGND.n1481 VGND.t520 17.4005
R5710 VGND.n1481 VGND.t135 17.4005
R5711 VGND.n1461 VGND.t44 17.4005
R5712 VGND.n1461 VGND.t339 17.4005
R5713 VGND.n1462 VGND.t341 17.4005
R5714 VGND.n1462 VGND.t362 17.4005
R5715 VGND.n1463 VGND.t247 17.4005
R5716 VGND.n1463 VGND.t353 17.4005
R5717 VGND.n1472 VGND.t351 17.4005
R5718 VGND.n1472 VGND.t197 17.4005
R5719 VGND.n1156 VGND.t530 17.4005
R5720 VGND.n1156 VGND.t76 17.4005
R5721 VGND.n1153 VGND.t210 17.4005
R5722 VGND.n1153 VGND.t208 17.4005
R5723 VGND.n1152 VGND.t167 17.4005
R5724 VGND.n1152 VGND.t499 17.4005
R5725 VGND.n1151 VGND.t334 17.4005
R5726 VGND.n1151 VGND.t151 17.4005
R5727 VGND.n1144 VGND.t289 17.4005
R5728 VGND.n1144 VGND.t420 17.4005
R5729 VGND.n1143 VGND.t418 17.4005
R5730 VGND.n1143 VGND.t291 17.4005
R5731 VGND.n1142 VGND.t295 17.4005
R5732 VGND.n1142 VGND.t458 17.4005
R5733 VGND.n1141 VGND.t147 17.4005
R5734 VGND.n1141 VGND.t490 17.4005
R5735 VGND.n1762 VGND.t234 17.1575
R5736 VGND.n241 VGND.t546 16.6727
R5737 VGND.n1024 VGND.t229 16.5844
R5738 VGND.t183 VGND.n1040 16.5844
R5739 VGND.n1830 VGND.t236 15.9478
R5740 VGND.n1728 VGND.n1727 15.3952
R5741 VGND.n1727 VGND.n1726 15.3952
R5742 VGND.n1303 VGND.n525 15.3952
R5743 VGND.n1726 VGND.n525 15.3952
R5744 VGND.n1328 VGND.n523 15.3952
R5745 VGND.n1726 VGND.n523 15.3952
R5746 VGND.n1353 VGND.n526 15.3952
R5747 VGND.n1726 VGND.n526 15.3952
R5748 VGND.n1378 VGND.n522 15.3952
R5749 VGND.n1726 VGND.n522 15.3952
R5750 VGND.n1223 VGND.n527 15.3952
R5751 VGND.n1726 VGND.n527 15.3952
R5752 VGND.n1260 VGND.n521 15.3952
R5753 VGND.n1726 VGND.n521 15.3952
R5754 VGND.n1725 VGND.n1724 15.3952
R5755 VGND.n1726 VGND.n1725 15.3952
R5756 VGND.n976 VGND.n781 15.2658
R5757 VGND.t141 VGND.n11 14.0522
R5758 VGND.n1754 VGND.n160 11.8985
R5759 VGND.t193 VGND.n588 11.842
R5760 VGND.t72 VGND.n612 11.842
R5761 VGND.t306 VGND.n636 11.842
R5762 VGND.t508 VGND.n660 11.842
R5763 VGND.t71 VGND.n684 11.842
R5764 VGND.n1069 VGND.t238 11.842
R5765 VGND.n1130 VGND.t474 11.0862
R5766 VGND.n1130 VGND.t84 11.0862
R5767 VGND.n1117 VGND.t22 11.0862
R5768 VGND.n1117 VGND.t185 11.0862
R5769 VGND.n1104 VGND.t173 11.0862
R5770 VGND.n1104 VGND.t144 11.0862
R5771 VGND.n1091 VGND.t239 11.0862
R5772 VGND.n1091 VGND.t179 11.0862
R5773 VGND.n1078 VGND.t293 11.0862
R5774 VGND.n1078 VGND.t45 11.0862
R5775 VGND.n720 VGND.t349 11.0862
R5776 VGND.n720 VGND.t113 11.0862
R5777 VGND.n1394 VGND.t21 10.6561
R5778 VGND.n588 VGND.t542 10.3303
R5779 VGND.n612 VGND.t336 10.3303
R5780 VGND.n636 VGND.t82 10.3303
R5781 VGND.n660 VGND.t433 10.3303
R5782 VGND.n684 VGND.t148 10.3303
R5783 VGND.t232 VGND.n1069 10.3303
R5784 VGND.n1020 VGND.n1019 8.89919
R5785 VGND.n1051 VGND.n1028 8.89919
R5786 VGND.n1041 VGND.n1036 8.89919
R5787 VGND.n1745 VGND.n332 8.89919
R5788 VGND.n990 VGND.t2 7.40866
R5789 VGND.n771 VGND.t478 6.73519
R5790 VGND.n1771 VGND 6.60769
R5791 VGND.n1747 VGND.n137 6.22424
R5792 VGND.n1748 VGND.n1747 6.06172
R5793 VGND.n1732 VGND.n513 5.90952
R5794 VGND.n515 VGND.t161 5.8005
R5795 VGND.n515 VGND.t251 5.8005
R5796 VGND.n1280 VGND.t301 5.8005
R5797 VGND.n1280 VGND.t92 5.8005
R5798 VGND.n1279 VGND.t452 5.8005
R5799 VGND.n1279 VGND.t165 5.8005
R5800 VGND.n1278 VGND.t317 5.8005
R5801 VGND.n1278 VGND.t129 5.8005
R5802 VGND.n1276 VGND.t219 5.8005
R5803 VGND.n1276 VGND.t95 5.8005
R5804 VGND.n1275 VGND.t194 5.8005
R5805 VGND.n1275 VGND.t157 5.8005
R5806 VGND.n1273 VGND.t162 5.8005
R5807 VGND.n1273 VGND.t94 5.8005
R5808 VGND.n1272 VGND.t195 5.8005
R5809 VGND.n1272 VGND.t160 5.8005
R5810 VGND.n1270 VGND.t91 5.8005
R5811 VGND.n1270 VGND.t335 5.8005
R5812 VGND.n1269 VGND.t425 5.8005
R5813 VGND.n1269 VGND.t93 5.8005
R5814 VGND.n1224 VGND.t471 5.8005
R5815 VGND.n1224 VGND.t218 5.8005
R5816 VGND.n1225 VGND.t217 5.8005
R5817 VGND.n1225 VGND.t168 5.8005
R5818 VGND.n1238 VGND.t155 5.8005
R5819 VGND.n1238 VGND.t470 5.8005
R5820 VGND.n1255 VGND.t96 5.8005
R5821 VGND.n1255 VGND.t254 5.8005
R5822 VGND.n569 VGND.t159 5.8005
R5823 VGND.n569 VGND.t451 5.8005
R5824 VGND.n568 VGND.t427 5.8005
R5825 VGND.n568 VGND.t99 5.8005
R5826 VGND.n582 VGND.n564 5.54333
R5827 VGND.n1129 VGND.n592 5.54333
R5828 VGND.n608 VGND.n607 5.54333
R5829 VGND.n1116 VGND.n616 5.54333
R5830 VGND.n632 VGND.n631 5.54333
R5831 VGND.n1103 VGND.n640 5.54333
R5832 VGND.n656 VGND.n655 5.54333
R5833 VGND.n1090 VGND.n664 5.54333
R5834 VGND.n680 VGND.n679 5.54333
R5835 VGND.n1077 VGND.n688 5.54333
R5836 VGND.n1070 VGND.n698 5.54333
R5837 VGND.n725 VGND.n715 5.54333
R5838 VGND.t21 VGND.n1168 5.45827
R5839 VGND.n990 VGND.t88 5.16377
R5840 VGND VGND.n1771 4.64147
R5841 VGND.n1769 VGND.n1768 4.6393
R5842 VGND.n1139 VGND.n1138 3.89165
R5843 VGND.n1732 VGND.n1731 3.78262
R5844 VGND.t8 VGND.n137 3.70013
R5845 VGND VGND.n1802 3.50128
R5846 VGND.n295 VGND.n285 3.46248
R5847 VGND.n299 VGND.n298 3.46248
R5848 VGND.n291 VGND.n290 3.46248
R5849 VGND.n294 VGND.n286 3.46248
R5850 VGND.n276 VGND.n212 3.46248
R5851 VGND.n280 VGND.n279 3.46248
R5852 VGND.n272 VGND.n271 3.46248
R5853 VGND.n275 VGND.n213 3.46248
R5854 VGND.n243 VGND.n0 3.46248
R5855 VGND.n246 VGND.n235 3.46248
R5856 VGND.n149 VGND.n148 3.46248
R5857 VGND.n992 VGND.n741 3.46248
R5858 VGND.n995 VGND.n738 3.46248
R5859 VGND.n983 VGND.n765 3.46248
R5860 VGND.n987 VGND.n986 3.46248
R5861 VGND.n965 VGND.n964 3.46248
R5862 VGND.n968 VGND.n795 3.46248
R5863 VGND.n960 VGND.n959 3.46248
R5864 VGND.n963 VGND.n798 3.46248
R5865 VGND.n943 VGND.n942 3.46248
R5866 VGND.n946 VGND.n809 3.46248
R5867 VGND.n938 VGND.n937 3.46248
R5868 VGND.n941 VGND.n812 3.46248
R5869 VGND.n921 VGND.n920 3.46248
R5870 VGND.n924 VGND.n823 3.46248
R5871 VGND.n916 VGND.n915 3.46248
R5872 VGND.n919 VGND.n826 3.46248
R5873 VGND.n899 VGND.n898 3.46248
R5874 VGND.n902 VGND.n837 3.46248
R5875 VGND.n894 VGND.n893 3.46248
R5876 VGND.n897 VGND.n840 3.46248
R5877 VGND.n877 VGND.n876 3.46248
R5878 VGND.n880 VGND.n851 3.46248
R5879 VGND.n872 VGND.n871 3.46248
R5880 VGND.n875 VGND.n854 3.46248
R5881 VGND.n1774 VGND.n1772 3.46248
R5882 VGND.n127 VGND.n125 3.46248
R5883 VGND.n121 VGND.n119 3.46248
R5884 VGND.n115 VGND.n113 3.46248
R5885 VGND.n109 VGND.n107 3.46248
R5886 VGND.n103 VGND.n101 3.46248
R5887 VGND.n97 VGND.n95 3.46248
R5888 VGND.n91 VGND.n89 3.46248
R5889 VGND.n86 VGND.n68 3.46248
R5890 VGND.n1805 VGND.n1803 3.46248
R5891 VGND.n65 VGND.n63 3.46248
R5892 VGND.n59 VGND.n57 3.46248
R5893 VGND.n53 VGND.n51 3.46248
R5894 VGND.n47 VGND.n45 3.46248
R5895 VGND.n41 VGND.n39 3.46248
R5896 VGND.n35 VGND.n33 3.46248
R5897 VGND.n29 VGND.n27 3.46248
R5898 VGND.n23 VGND.n21 3.46248
R5899 VGND.n472 VGND.n471 3.46248
R5900 VGND.n469 VGND.n467 3.46248
R5901 VGND.n463 VGND.n461 3.46248
R5902 VGND.n457 VGND.n455 3.46248
R5903 VGND.n451 VGND.n449 3.46248
R5904 VGND.n445 VGND.n443 3.46248
R5905 VGND.n439 VGND.n437 3.46248
R5906 VGND.n433 VGND.n431 3.46248
R5907 VGND.n427 VGND.n425 3.46248
R5908 VGND.n421 VGND.n419 3.46248
R5909 VGND.n415 VGND.n413 3.46248
R5910 VGND.n409 VGND.n407 3.46248
R5911 VGND.n403 VGND.n401 3.46248
R5912 VGND.n397 VGND.n395 3.46248
R5913 VGND.n391 VGND.n389 3.46248
R5914 VGND.n385 VGND.n383 3.46248
R5915 VGND.n379 VGND.n377 3.46248
R5916 VGND.n374 VGND.n367 3.46248
R5917 VGND.n370 VGND.n369 3.46248
R5918 VGND.n513 VGND.n340 3.46248
R5919 VGND.n154 VGND.n153 3.46248
R5920 VGND.n1769 VGND.n4 3.07882
R5921 VGND.n1770 VGND.n1769 3.02279
R5922 VGND.n1706 VGND.n1705 3.0154
R5923 VGND.n1731 VGND 2.95362
R5924 VGND.n1750 VGND.n164 2.913
R5925 VGND.n1758 VGND.n1757 2.913
R5926 VGND.n257 VGND.n221 2.913
R5927 VGND.n253 VGND.n229 2.913
R5928 VGND.n323 VGND.n175 2.82278
R5929 VGND.n319 VGND.n181 2.82278
R5930 VGND.n322 VGND.n176 2.82278
R5931 VGND.n309 VGND.n195 2.82278
R5932 VGND.n289 VGND.n194 2.82278
R5933 VGND.n305 VGND.n203 2.82278
R5934 VGND.n308 VGND.n199 2.82278
R5935 VGND.n1011 VGND.n732 2.82278
R5936 VGND.n1007 VGND.n996 2.82278
R5937 VGND.n1010 VGND.n733 2.82278
R5938 VGND.n978 VGND.n769 2.82278
R5939 VGND.n982 VGND.n766 2.82278
R5940 VGND.n969 VGND.n794 2.82278
R5941 VGND.n973 VGND.n972 2.82278
R5942 VGND.n954 VGND.n952 2.82278
R5943 VGND.n958 VGND.n801 2.82278
R5944 VGND.n948 VGND.n947 2.82278
R5945 VGND.n951 VGND.n804 2.82278
R5946 VGND.n932 VGND.n930 2.82278
R5947 VGND.n936 VGND.n815 2.82278
R5948 VGND.n926 VGND.n925 2.82278
R5949 VGND.n929 VGND.n818 2.82278
R5950 VGND.n910 VGND.n908 2.82278
R5951 VGND.n914 VGND.n829 2.82278
R5952 VGND.n904 VGND.n903 2.82278
R5953 VGND.n907 VGND.n832 2.82278
R5954 VGND.n888 VGND.n886 2.82278
R5955 VGND.n892 VGND.n843 2.82278
R5956 VGND.n882 VGND.n881 2.82278
R5957 VGND.n885 VGND.n846 2.82278
R5958 VGND.n1015 VGND.n1014 2.82278
R5959 VGND.n327 VGND.n326 2.82278
R5960 VGND.n1801 VGND.n69 2.768
R5961 VGND.n1644 VGND.n74 2.768
R5962 VGND.n1658 VGND.n1645 2.768
R5963 VGND.n1663 VGND.n1634 2.768
R5964 VGND.n1664 VGND.n1633 2.768
R5965 VGND.n1671 VGND.n1670 2.768
R5966 VGND.n1676 VGND.n1618 2.768
R5967 VGND.n1681 VGND.n1610 2.768
R5968 VGND.n1682 VGND.n1609 2.768
R5969 VGND.n1689 VGND.n1688 2.768
R5970 VGND.n1694 VGND.n1594 2.768
R5971 VGND.n1699 VGND.n1586 2.768
R5972 VGND.n1700 VGND.n1585 2.768
R5973 VGND.n1531 VGND.n1530 2.768
R5974 VGND.n1542 VGND.n1523 2.768
R5975 VGND.n1544 VGND.n1543 2.768
R5976 VGND.n1517 VGND.n1411 2.768
R5977 VGND.n1516 VGND.n1412 2.768
R5978 VGND.n1511 VGND.n1510 2.768
R5979 VGND.n1507 VGND.n1424 2.768
R5980 VGND.n1502 VGND.n1501 2.768
R5981 VGND.n1498 VGND.n1436 2.768
R5982 VGND.n1493 VGND.n1492 2.768
R5983 VGND.n1489 VGND.n1448 2.768
R5984 VGND.n1484 VGND.n1483 2.768
R5985 VGND.n1480 VGND.n1460 2.768
R5986 VGND.n1475 VGND.n1474 2.768
R5987 VGND.n1552 VGND.n1158 2.768
R5988 VGND.n1557 VGND.n1150 2.768
R5989 VGND.n1558 VGND.n1149 2.768
R5990 VGND.n1565 VGND.n1564 2.768
R5991 VGND.n1407 VGND.n1401 2.52995
R5992 VGND.n1418 VGND.n1417 2.52995
R5993 VGND.n1430 VGND.n1429 2.52995
R5994 VGND.n1442 VGND.n1441 2.52995
R5995 VGND.n1454 VGND.n1453 2.52995
R5996 VGND.n1466 VGND.n1465 2.52995
R5997 VGND.n1159 VGND.n1155 2.52995
R5998 VGND.n1145 VGND.n566 2.52995
R5999 VGND.n1646 VGND.n1639 2.52995
R6000 VGND.n1647 VGND.n1627 2.52995
R6001 VGND.n1619 VGND.n1615 2.52995
R6002 VGND.n1620 VGND.n1603 2.52995
R6003 VGND.n1595 VGND.n1591 2.52995
R6004 VGND.n1596 VGND.n1579 2.52995
R6005 VGND.n1537 VGND.n1533 2.52995
R6006 VGND.n1796 VGND.n75 2.52995
R6007 VGND.n1731 VGND 2.40675
R6008 VGND.n1140 VGND.n1139 2.3961
R6009 VGND.n1752 VGND.n164 2.3255
R6010 VGND.n1757 VGND.n1756 2.3255
R6011 VGND.n1775 VGND.n128 2.3255
R6012 VGND.n1777 VGND.n122 2.3255
R6013 VGND.n1779 VGND.n116 2.3255
R6014 VGND.n1781 VGND.n110 2.3255
R6015 VGND.n1783 VGND.n104 2.3255
R6016 VGND.n1785 VGND.n98 2.3255
R6017 VGND.n1787 VGND.n92 2.3255
R6018 VGND.n1789 VGND.n87 2.3255
R6019 VGND.n1806 VGND.n66 2.3255
R6020 VGND.n1808 VGND.n60 2.3255
R6021 VGND.n1810 VGND.n54 2.3255
R6022 VGND.n1812 VGND.n48 2.3255
R6023 VGND.n1814 VGND.n42 2.3255
R6024 VGND.n1816 VGND.n36 2.3255
R6025 VGND.n1818 VGND.n30 2.3255
R6026 VGND.n1820 VGND.n24 2.3255
R6027 VGND.n1822 VGND.n19 2.3255
R6028 VGND.n475 VGND.n474 2.3255
R6029 VGND.n477 VGND.n464 2.3255
R6030 VGND.n479 VGND.n458 2.3255
R6031 VGND.n481 VGND.n452 2.3255
R6032 VGND.n483 VGND.n446 2.3255
R6033 VGND.n485 VGND.n440 2.3255
R6034 VGND.n487 VGND.n434 2.3255
R6035 VGND.n489 VGND.n428 2.3255
R6036 VGND.n491 VGND.n422 2.3255
R6037 VGND.n493 VGND.n416 2.3255
R6038 VGND.n495 VGND.n410 2.3255
R6039 VGND.n497 VGND.n404 2.3255
R6040 VGND.n499 VGND.n398 2.3255
R6041 VGND.n501 VGND.n392 2.3255
R6042 VGND.n503 VGND.n386 2.3255
R6043 VGND.n505 VGND.n380 2.3255
R6044 VGND.n507 VGND.n375 2.3255
R6045 VGND.n372 VGND.n371 2.3255
R6046 VGND.n512 VGND.n511 2.3255
R6047 VGND.n265 VGND.n221 2.3255
R6048 VGND.n231 VGND.n229 2.3255
R6049 VGND.n985 VGND.n764 2.3255
R6050 VGND.n994 VGND.n993 2.3255
R6051 VGND.n962 VGND.n961 2.3255
R6052 VGND.n967 VGND.n966 2.3255
R6053 VGND.n940 VGND.n939 2.3255
R6054 VGND.n945 VGND.n944 2.3255
R6055 VGND.n918 VGND.n917 2.3255
R6056 VGND.n923 VGND.n922 2.3255
R6057 VGND.n896 VGND.n895 2.3255
R6058 VGND.n901 VGND.n900 2.3255
R6059 VGND.n874 VGND.n873 2.3255
R6060 VGND.n879 VGND.n878 2.3255
R6061 VGND.n144 VGND.n143 2.3255
R6062 VGND.n293 VGND.n292 2.3255
R6063 VGND.n297 VGND.n284 2.3255
R6064 VGND.n274 VGND.n273 2.3255
R6065 VGND.n278 VGND.n211 2.3255
R6066 VGND.n245 VGND.n244 2.3255
R6067 VGND.n1139 VGND.n573 2.28621
R6068 VGND.n239 VGND.n238 2.17513
R6069 VGND.n1832 VGND.n4 2.15467
R6070 VGND.n1768 VGND.n130 2.15467
R6071 VGND.n1835 VGND.n1 2.1305
R6072 VGND.n132 VGND.n131 2.1305
R6073 VGND.n1712 VGND.n537 2.07965
R6074 VGND.n869 VGND.n858 1.95084
R6075 VGND.n865 VGND.n141 1.95084
R6076 VGND.n269 VGND.n216 1.95084
R6077 VGND.n251 VGND.n250 1.95084
R6078 VGND.n1766 VGND.n1765 1.8605
R6079 VGND.n1834 VGND.n1833 1.8605
R6080 VGND.n1730 VGND.n514 1.56378
R6081 VGND.n1302 VGND.n1284 1.56378
R6082 VGND.n1327 VGND.n1309 1.56378
R6083 VGND.n1352 VGND.n1334 1.56378
R6084 VGND.n1377 VGND.n1359 1.56378
R6085 VGND.n1387 VGND.n1384 1.56378
R6086 VGND.n1262 VGND.n1237 1.56378
R6087 VGND.n1723 VGND.n532 1.56378
R6088 VGND.n270 VGND.n269 1.52133
R6089 VGND VGND.n1557 1.3768
R6090 VGND.n1474 VGND 1.3768
R6091 VGND.n1483 VGND 1.3768
R6092 VGND.n1492 VGND 1.3768
R6093 VGND.n1501 VGND 1.3768
R6094 VGND.n1510 VGND 1.3768
R6095 VGND.n1517 VGND 1.3768
R6096 VGND VGND.n1542 1.3768
R6097 VGND.n1283 VGND.n517 1.37182
R6098 VGND.n1308 VGND.n1277 1.37182
R6099 VGND.n1333 VGND.n1274 1.37182
R6100 VGND.n1358 VGND.n1271 1.37182
R6101 VGND.n1383 VGND.n1268 1.37182
R6102 VGND.n1263 VGND.n1234 1.37182
R6103 VGND.n1259 VGND.n1258 1.37182
R6104 VGND.n573 VGND.n530 1.37182
R6105 VGND.n1009 VGND.n1008 1.32907
R6106 VGND.n1012 VGND.n727 1.32907
R6107 VGND.n971 VGND.n791 1.32907
R6108 VGND.n980 VGND.n979 1.32907
R6109 VGND.n950 VGND.n949 1.32907
R6110 VGND.n956 VGND.n955 1.32907
R6111 VGND.n928 VGND.n927 1.32907
R6112 VGND.n934 VGND.n933 1.32907
R6113 VGND.n906 VGND.n905 1.32907
R6114 VGND.n912 VGND.n911 1.32907
R6115 VGND.n884 VGND.n883 1.32907
R6116 VGND.n890 VGND.n889 1.32907
R6117 VGND.n321 VGND.n320 1.32907
R6118 VGND.n324 VGND.n170 1.32907
R6119 VGND.n307 VGND.n306 1.32907
R6120 VGND.n311 VGND.n310 1.32907
R6121 VGND.n870 VGND.n869 1.30085
R6122 VGND.n1140 VGND 1.21891
R6123 VGND.n1014 VGND.n729 0.959726
R6124 VGND.n326 VGND.n172 0.959726
R6125 VGND.n249 VGND.n234 0.957022
R6126 VGND.n268 VGND.n218 0.957022
R6127 VGND.n864 VGND.n862 0.957022
R6128 VGND.n868 VGND.n860 0.957022
R6129 VGND.n532 VGND.n531 0.785098
R6130 VGND.n1262 VGND.n1261 0.785098
R6131 VGND.n1384 VGND.n1267 0.785098
R6132 VGND.n1379 VGND.n1359 0.785098
R6133 VGND.n1354 VGND.n1334 0.785098
R6134 VGND.n1329 VGND.n1309 0.785098
R6135 VGND.n1304 VGND.n1284 0.785098
R6136 VGND.n1730 VGND.n1729 0.785098
R6137 VGND.n1771 VGND.n1770 0.738047
R6138 VGND.n202 VGND.n201 0.685283
R6139 VGND.n198 VGND.n197 0.685283
R6140 VGND.n179 VGND.n178 0.685283
R6141 VGND.n325 VGND.n174 0.685283
R6142 VGND.n849 VGND.n848 0.685283
R6143 VGND.n891 VGND.n845 0.685283
R6144 VGND.n835 VGND.n834 0.685283
R6145 VGND.n913 VGND.n831 0.685283
R6146 VGND.n821 VGND.n820 0.685283
R6147 VGND.n935 VGND.n817 0.685283
R6148 VGND.n807 VGND.n806 0.685283
R6149 VGND.n957 VGND.n803 0.685283
R6150 VGND.n970 VGND.n793 0.685283
R6151 VGND.n981 VGND.n768 0.685283
R6152 VGND.n736 VGND.n735 0.685283
R6153 VGND.n1013 VGND.n731 0.685283
R6154 VGND VGND.n1125 0.669618
R6155 VGND VGND.n1112 0.669618
R6156 VGND VGND.n1099 0.669618
R6157 VGND VGND.n1086 0.669618
R6158 VGND VGND.n1073 0.669618
R6159 VGND VGND.n1060 0.669618
R6160 VGND VGND.n1047 0.669618
R6161 VGND.n1798 VGND.n1797 0.58175
R6162 VGND.n1660 VGND.n1659 0.58175
R6163 VGND.n1667 VGND.n1628 0.58175
R6164 VGND.n1678 VGND.n1677 0.58175
R6165 VGND.n1685 VGND.n1604 0.58175
R6166 VGND.n1696 VGND.n1695 0.58175
R6167 VGND.n1703 VGND.n1580 0.58175
R6168 VGND.n1539 VGND.n1538 0.58175
R6169 VGND.n1520 VGND.n1402 0.58175
R6170 VGND.n1513 VGND.n1512 0.58175
R6171 VGND.n1504 VGND.n1503 0.58175
R6172 VGND.n1495 VGND.n1494 0.58175
R6173 VGND.n1486 VGND.n1485 0.58175
R6174 VGND.n1477 VGND.n1476 0.58175
R6175 VGND.n1554 VGND.n1553 0.58175
R6176 VGND.n1561 VGND.n567 0.58175
R6177 VGND.n1037 VGND.n338 0.58175
R6178 VGND.n1057 VGND.n1056 0.58175
R6179 VGND.n1083 VGND.n1082 0.58175
R6180 VGND.n1096 VGND.n1095 0.58175
R6181 VGND.n1109 VGND.n1108 0.58175
R6182 VGND.n1122 VGND.n1121 0.58175
R6183 VGND.n1135 VGND.n1134 0.58175
R6184 VGND.n1066 VGND.n1065 0.58175
R6185 VGND.n729 VGND 0.578086
R6186 VGND.n172 VGND 0.578086
R6187 VGND.n1564 VGND.n1140 0.53826
R6188 VGND VGND.n154 0.523938
R6189 VGND VGND.n246 0.523938
R6190 VGND VGND.n532 0.522821
R6191 VGND VGND.n1262 0.522821
R6192 VGND.n1384 VGND 0.522821
R6193 VGND.n1359 VGND 0.522821
R6194 VGND.n1334 VGND 0.522821
R6195 VGND.n1309 VGND 0.522821
R6196 VGND.n1284 VGND 0.522821
R6197 VGND VGND.n1730 0.522821
R6198 VGND.n1729 VGND.n1728 0.517167
R6199 VGND.n1304 VGND.n1303 0.517167
R6200 VGND.n1329 VGND.n1328 0.517167
R6201 VGND.n1354 VGND.n1353 0.517167
R6202 VGND.n1379 VGND.n1378 0.517167
R6203 VGND.n1267 VGND.n1223 0.517167
R6204 VGND.n1261 VGND.n1260 0.517167
R6205 VGND.n1724 VGND.n531 0.517167
R6206 VGND.n983 VGND 0.479667
R6207 VGND.n959 VGND 0.479667
R6208 VGND.n937 VGND 0.479667
R6209 VGND.n915 VGND 0.479667
R6210 VGND.n893 VGND 0.479667
R6211 VGND.n290 VGND 0.479667
R6212 VGND VGND.n995 0.466646
R6213 VGND VGND.n968 0.466646
R6214 VGND VGND.n946 0.466646
R6215 VGND VGND.n924 0.466646
R6216 VGND VGND.n902 0.466646
R6217 VGND VGND.n880 0.466646
R6218 VGND.n298 VGND 0.466646
R6219 VGND.n279 VGND 0.466646
R6220 VGND.n148 VGND 0.463123
R6221 VGND VGND.n0 0.463123
R6222 VGND.n1258 VGND 0.455857
R6223 VGND.n1263 VGND 0.455857
R6224 VGND VGND.n1383 0.455857
R6225 VGND VGND.n1358 0.455857
R6226 VGND VGND.n1333 0.455857
R6227 VGND VGND.n1308 0.455857
R6228 VGND VGND.n1283 0.455857
R6229 VGND.n866 VGND.n164 0.440404
R6230 VGND.n1757 VGND.n155 0.440404
R6231 VGND.n221 VGND.n219 0.440404
R6232 VGND.n247 VGND.n229 0.440404
R6233 VGND.n1011 VGND.n1010 0.430188
R6234 VGND.n972 VGND.n769 0.430188
R6235 VGND.n952 VGND.n951 0.430188
R6236 VGND.n930 VGND.n929 0.430188
R6237 VGND.n908 VGND.n907 0.430188
R6238 VGND.n886 VGND.n885 0.430188
R6239 VGND.n323 VGND.n322 0.430188
R6240 VGND.n309 VGND.n308 0.430188
R6241 VGND.n1802 VGND 0.426281
R6242 VGND.n863 VGND.n156 0.423227
R6243 VGND.n867 VGND.n163 0.423227
R6244 VGND.n248 VGND.n232 0.423227
R6245 VGND.n267 VGND.n266 0.423227
R6246 VGND.n271 VGND.n270 0.383313
R6247 VGND.n1037 VGND.n336 0.376971
R6248 VGND.n1056 VGND.n1055 0.376971
R6249 VGND.n1082 VGND.n1081 0.376971
R6250 VGND.n1095 VGND.n1094 0.376971
R6251 VGND.n1108 VGND.n1107 0.376971
R6252 VGND.n1121 VGND.n1120 0.376971
R6253 VGND.n1134 VGND.n1133 0.376971
R6254 VGND.n1066 VGND.n700 0.376971
R6255 VGND.n1012 VGND.n1011 0.359875
R6256 VGND.n1010 VGND.n1009 0.359875
R6257 VGND.n980 VGND.n769 0.359875
R6258 VGND.n972 VGND.n971 0.359875
R6259 VGND.n956 VGND.n952 0.359875
R6260 VGND.n951 VGND.n950 0.359875
R6261 VGND.n934 VGND.n930 0.359875
R6262 VGND.n929 VGND.n928 0.359875
R6263 VGND.n912 VGND.n908 0.359875
R6264 VGND.n907 VGND.n906 0.359875
R6265 VGND.n890 VGND.n886 0.359875
R6266 VGND.n885 VGND.n884 0.359875
R6267 VGND.n324 VGND.n323 0.359875
R6268 VGND.n322 VGND.n321 0.359875
R6269 VGND.n310 VGND.n309 0.359875
R6270 VGND.n308 VGND.n307 0.359875
R6271 VGND.n1137 VGND.n1136 0.324029
R6272 VGND.n595 VGND.n594 0.324029
R6273 VGND.n1124 VGND.n1123 0.324029
R6274 VGND.n619 VGND.n618 0.324029
R6275 VGND.n1111 VGND.n1110 0.324029
R6276 VGND.n643 VGND.n642 0.324029
R6277 VGND.n1098 VGND.n1097 0.324029
R6278 VGND.n667 VGND.n666 0.324029
R6279 VGND.n1085 VGND.n1084 0.324029
R6280 VGND.n691 VGND.n690 0.324029
R6281 VGND.n701 VGND.n693 0.324029
R6282 VGND.n1063 VGND.n1062 0.324029
R6283 VGND.n1059 VGND.n1058 0.324029
R6284 VGND.n1031 VGND.n1030 0.324029
R6285 VGND.n1046 VGND.n1045 0.324029
R6286 VGND.n1735 VGND.n1734 0.324029
R6287 VGND.n871 VGND.n870 0.323417
R6288 VGND.n866 VGND 0.306056
R6289 VGND.n155 VGND 0.306056
R6290 VGND VGND.n219 0.306056
R6291 VGND.n247 VGND 0.306056
R6292 VGND.n1770 VGND 0.284263
R6293 VGND.n1704 VGND.n1703 0.247896
R6294 VGND.n1703 VGND.n1702 0.247896
R6295 VGND.n1701 VGND.n1700 0.247896
R6296 VGND.n1699 VGND.n1698 0.247896
R6297 VGND.n1697 VGND.n1696 0.247896
R6298 VGND.n1696 VGND.n1590 0.247896
R6299 VGND.n1594 VGND.n1593 0.247896
R6300 VGND.n1688 VGND.n1687 0.247896
R6301 VGND.n1686 VGND.n1685 0.247896
R6302 VGND.n1685 VGND.n1684 0.247896
R6303 VGND.n1683 VGND.n1682 0.247896
R6304 VGND.n1681 VGND.n1680 0.247896
R6305 VGND.n1679 VGND.n1678 0.247896
R6306 VGND.n1678 VGND.n1614 0.247896
R6307 VGND.n1618 VGND.n1617 0.247896
R6308 VGND.n1670 VGND.n1669 0.247896
R6309 VGND.n1668 VGND.n1667 0.247896
R6310 VGND.n1667 VGND.n1666 0.247896
R6311 VGND.n1665 VGND.n1664 0.247896
R6312 VGND.n1663 VGND.n1662 0.247896
R6313 VGND.n1661 VGND.n1660 0.247896
R6314 VGND.n1660 VGND.n1638 0.247896
R6315 VGND.n1645 VGND.n1641 0.247896
R6316 VGND.n1644 VGND.n1643 0.247896
R6317 VGND.n1798 VGND.n73 0.247896
R6318 VGND.n1799 VGND.n1798 0.247896
R6319 VGND.n1801 VGND.n1800 0.247896
R6320 VGND.n1564 VGND.n1563 0.247896
R6321 VGND.n1562 VGND.n1561 0.247896
R6322 VGND.n1561 VGND.n1560 0.247896
R6323 VGND.n1559 VGND.n1558 0.247896
R6324 VGND.n1557 VGND.n1556 0.247896
R6325 VGND.n1555 VGND.n1554 0.247896
R6326 VGND.n1554 VGND.n1154 0.247896
R6327 VGND.n1158 VGND.n1157 0.247896
R6328 VGND.n1474 VGND.n1473 0.247896
R6329 VGND.n1477 VGND.n1464 0.247896
R6330 VGND.n1478 VGND.n1477 0.247896
R6331 VGND.n1480 VGND.n1479 0.247896
R6332 VGND.n1483 VGND.n1482 0.247896
R6333 VGND.n1486 VGND.n1452 0.247896
R6334 VGND.n1487 VGND.n1486 0.247896
R6335 VGND.n1489 VGND.n1488 0.247896
R6336 VGND.n1492 VGND.n1491 0.247896
R6337 VGND.n1495 VGND.n1440 0.247896
R6338 VGND.n1496 VGND.n1495 0.247896
R6339 VGND.n1498 VGND.n1497 0.247896
R6340 VGND.n1501 VGND.n1500 0.247896
R6341 VGND.n1504 VGND.n1428 0.247896
R6342 VGND.n1505 VGND.n1504 0.247896
R6343 VGND.n1507 VGND.n1506 0.247896
R6344 VGND.n1510 VGND.n1509 0.247896
R6345 VGND.n1513 VGND.n1416 0.247896
R6346 VGND.n1514 VGND.n1513 0.247896
R6347 VGND.n1516 VGND.n1515 0.247896
R6348 VGND.n1518 VGND.n1517 0.247896
R6349 VGND.n1520 VGND.n1519 0.247896
R6350 VGND.n1521 VGND.n1520 0.247896
R6351 VGND.n1543 VGND.n1522 0.247896
R6352 VGND.n1542 VGND.n1541 0.247896
R6353 VGND.n1540 VGND.n1539 0.247896
R6354 VGND.n1539 VGND.n1527 0.247896
R6355 VGND.n1530 VGND.n1529 0.247896
R6356 VGND.n570 VGND.n531 0.246036
R6357 VGND.n1261 VGND.n1239 0.246036
R6358 VGND.n1267 VGND.n1266 0.246036
R6359 VGND.n1380 VGND.n1379 0.246036
R6360 VGND.n1355 VGND.n1354 0.246036
R6361 VGND.n1330 VGND.n1329 0.246036
R6362 VGND.n1305 VGND.n1304 0.246036
R6363 VGND.n1729 VGND.n516 0.246036
R6364 VGND.n1138 VGND.n1137 0.239471
R6365 VGND.n1125 VGND.n1124 0.239471
R6366 VGND.n1112 VGND.n1111 0.239471
R6367 VGND.n1099 VGND.n1098 0.239471
R6368 VGND.n1086 VGND.n1085 0.239471
R6369 VGND.n1073 VGND.n693 0.239471
R6370 VGND.n1060 VGND.n1059 0.239471
R6371 VGND.n1047 VGND.n1046 0.239471
R6372 VGND.n1126 VGND.n595 0.232118
R6373 VGND.n1113 VGND.n619 0.232118
R6374 VGND.n1100 VGND.n643 0.232118
R6375 VGND.n1087 VGND.n667 0.232118
R6376 VGND.n1074 VGND.n691 0.232118
R6377 VGND.n1062 VGND.n1061 0.232118
R6378 VGND.n1048 VGND.n1031 0.232118
R6379 VGND.n1734 VGND.n1733 0.232118
R6380 VGND.n1766 VGND.n131 0.230892
R6381 VGND.n1835 VGND.n1834 0.230892
R6382 VGND.n1705 VGND.n1704 0.229667
R6383 VGND.n1702 VGND.n1701 0.229667
R6384 VGND.n1698 VGND.n1697 0.229667
R6385 VGND.n1593 VGND.n1590 0.229667
R6386 VGND.n1687 VGND.n1686 0.229667
R6387 VGND.n1684 VGND.n1683 0.229667
R6388 VGND.n1680 VGND.n1679 0.229667
R6389 VGND.n1617 VGND.n1614 0.229667
R6390 VGND.n1669 VGND.n1668 0.229667
R6391 VGND.n1666 VGND.n1665 0.229667
R6392 VGND.n1662 VGND.n1661 0.229667
R6393 VGND.n1641 VGND.n1638 0.229667
R6394 VGND.n1643 VGND.n73 0.229667
R6395 VGND.n1800 VGND.n1799 0.229667
R6396 VGND.n1563 VGND.n1562 0.229667
R6397 VGND.n1560 VGND.n1559 0.229667
R6398 VGND.n1556 VGND.n1555 0.229667
R6399 VGND.n1157 VGND.n1154 0.229667
R6400 VGND.n1473 VGND.n1464 0.229667
R6401 VGND.n1479 VGND.n1478 0.229667
R6402 VGND.n1482 VGND.n1452 0.229667
R6403 VGND.n1488 VGND.n1487 0.229667
R6404 VGND.n1491 VGND.n1440 0.229667
R6405 VGND.n1497 VGND.n1496 0.229667
R6406 VGND.n1500 VGND.n1428 0.229667
R6407 VGND.n1506 VGND.n1505 0.229667
R6408 VGND.n1509 VGND.n1416 0.229667
R6409 VGND.n1515 VGND.n1514 0.229667
R6410 VGND.n1519 VGND.n1518 0.229667
R6411 VGND.n1522 VGND.n1521 0.229667
R6412 VGND.n1541 VGND.n1540 0.229667
R6413 VGND.n1529 VGND.n1527 0.229667
R6414 VGND.n1013 VGND.n1012 0.229667
R6415 VGND.n1009 VGND.n736 0.229667
R6416 VGND.n981 VGND.n980 0.229667
R6417 VGND.n971 VGND.n970 0.229667
R6418 VGND.n957 VGND.n956 0.229667
R6419 VGND.n950 VGND.n807 0.229667
R6420 VGND.n935 VGND.n934 0.229667
R6421 VGND.n928 VGND.n821 0.229667
R6422 VGND.n913 VGND.n912 0.229667
R6423 VGND.n906 VGND.n835 0.229667
R6424 VGND.n891 VGND.n890 0.229667
R6425 VGND.n884 VGND.n849 0.229667
R6426 VGND.n325 VGND.n324 0.229667
R6427 VGND.n321 VGND.n179 0.229667
R6428 VGND.n310 VGND.n198 0.229667
R6429 VGND.n307 VGND.n202 0.229667
R6430 VGND.n781 VGND.t2 0.22499
R6431 VGND.n1802 VGND.n68 0.212219
R6432 VGND.n572 VGND.n571 0.196929
R6433 VGND.n571 VGND.n570 0.196929
R6434 VGND.n1257 VGND.n1256 0.196929
R6435 VGND.n1256 VGND.n1239 0.196929
R6436 VGND.n1265 VGND.n1264 0.196929
R6437 VGND.n1266 VGND.n1265 0.196929
R6438 VGND.n1382 VGND.n1381 0.196929
R6439 VGND.n1381 VGND.n1380 0.196929
R6440 VGND.n1357 VGND.n1356 0.196929
R6441 VGND.n1356 VGND.n1355 0.196929
R6442 VGND.n1332 VGND.n1331 0.196929
R6443 VGND.n1331 VGND.n1330 0.196929
R6444 VGND.n1307 VGND.n1306 0.196929
R6445 VGND.n1306 VGND.n1305 0.196929
R6446 VGND.n1282 VGND.n1281 0.196929
R6447 VGND.n1281 VGND.n516 0.196929
R6448 VGND VGND.n982 0.191906
R6449 VGND VGND.n958 0.191906
R6450 VGND VGND.n936 0.191906
R6451 VGND VGND.n914 0.191906
R6452 VGND VGND.n892 0.191906
R6453 VGND VGND.n289 0.191906
R6454 VGND.n87 VGND.n68 0.189302
R6455 VGND.n92 VGND.n91 0.189302
R6456 VGND.n98 VGND.n97 0.189302
R6457 VGND.n104 VGND.n103 0.189302
R6458 VGND.n110 VGND.n109 0.189302
R6459 VGND.n116 VGND.n115 0.189302
R6460 VGND.n122 VGND.n121 0.189302
R6461 VGND.n128 VGND.n127 0.189302
R6462 VGND.n513 VGND.n512 0.189302
R6463 VGND.n372 VGND.n370 0.189302
R6464 VGND.n375 VGND.n374 0.189302
R6465 VGND.n380 VGND.n379 0.189302
R6466 VGND.n386 VGND.n385 0.189302
R6467 VGND.n392 VGND.n391 0.189302
R6468 VGND.n398 VGND.n397 0.189302
R6469 VGND.n404 VGND.n403 0.189302
R6470 VGND.n410 VGND.n409 0.189302
R6471 VGND.n416 VGND.n415 0.189302
R6472 VGND.n422 VGND.n421 0.189302
R6473 VGND.n428 VGND.n427 0.189302
R6474 VGND.n434 VGND.n433 0.189302
R6475 VGND.n440 VGND.n439 0.189302
R6476 VGND.n446 VGND.n445 0.189302
R6477 VGND.n452 VGND.n451 0.189302
R6478 VGND.n458 VGND.n457 0.189302
R6479 VGND.n464 VGND.n463 0.189302
R6480 VGND.n474 VGND.n469 0.189302
R6481 VGND.n472 VGND.n19 0.189302
R6482 VGND.n24 VGND.n23 0.189302
R6483 VGND.n30 VGND.n29 0.189302
R6484 VGND.n36 VGND.n35 0.189302
R6485 VGND.n42 VGND.n41 0.189302
R6486 VGND.n48 VGND.n47 0.189302
R6487 VGND.n54 VGND.n53 0.189302
R6488 VGND.n60 VGND.n59 0.189302
R6489 VGND.n66 VGND.n65 0.189302
R6490 VGND.n995 VGND.n994 0.189302
R6491 VGND.n986 VGND.n985 0.189302
R6492 VGND.n968 VGND.n967 0.189302
R6493 VGND.n963 VGND.n962 0.189302
R6494 VGND.n946 VGND.n945 0.189302
R6495 VGND.n941 VGND.n940 0.189302
R6496 VGND.n924 VGND.n923 0.189302
R6497 VGND.n919 VGND.n918 0.189302
R6498 VGND.n902 VGND.n901 0.189302
R6499 VGND.n897 VGND.n896 0.189302
R6500 VGND.n880 VGND.n879 0.189302
R6501 VGND.n875 VGND.n874 0.189302
R6502 VGND.n154 VGND.n143 0.189302
R6503 VGND.n298 VGND.n297 0.189302
R6504 VGND.n294 VGND.n293 0.189302
R6505 VGND.n279 VGND.n278 0.189302
R6506 VGND.n275 VGND.n274 0.189302
R6507 VGND.n246 VGND.n245 0.189302
R6508 VGND VGND.n1732 0.172069
R6509 VGND.n869 VGND.n868 0.169771
R6510 VGND.n865 VGND.n864 0.169771
R6511 VGND.n269 VGND.n268 0.169771
R6512 VGND.n250 VGND.n249 0.169771
R6513 VGND.n868 VGND.n867 0.168035
R6514 VGND.n864 VGND.n863 0.168035
R6515 VGND.n268 VGND.n267 0.168035
R6516 VGND.n249 VGND.n248 0.168035
R6517 VGND VGND.n865 0.15675
R6518 VGND.n250 VGND 0.15675
R6519 VGND.n1700 VGND 0.147635
R6520 VGND VGND.n1594 0.147635
R6521 VGND.n1682 VGND 0.147635
R6522 VGND VGND.n1618 0.147635
R6523 VGND.n1664 VGND 0.147635
R6524 VGND.n1645 VGND 0.147635
R6525 VGND VGND.n1801 0.147635
R6526 VGND.n1558 VGND 0.147635
R6527 VGND VGND.n1158 0.147635
R6528 VGND VGND.n1480 0.147635
R6529 VGND VGND.n1489 0.147635
R6530 VGND VGND.n1498 0.147635
R6531 VGND VGND.n1507 0.147635
R6532 VGND VGND.n1516 0.147635
R6533 VGND.n1543 VGND 0.147635
R6534 VGND.n1530 VGND 0.147635
R6535 VGND.n573 VGND.n572 0.146705
R6536 VGND.n1258 VGND.n1257 0.146705
R6537 VGND.n1264 VGND.n1263 0.146705
R6538 VGND.n1383 VGND.n1382 0.146705
R6539 VGND.n1358 VGND.n1357 0.146705
R6540 VGND.n1333 VGND.n1332 0.146705
R6541 VGND.n1308 VGND.n1307 0.146705
R6542 VGND.n1283 VGND.n1282 0.146705
R6543 VGND.n986 VGND.n741 0.141125
R6544 VGND.n964 VGND.n963 0.141125
R6545 VGND.n942 VGND.n941 0.141125
R6546 VGND.n920 VGND.n919 0.141125
R6547 VGND.n898 VGND.n897 0.141125
R6548 VGND.n876 VGND.n875 0.141125
R6549 VGND.n295 VGND.n294 0.141125
R6550 VGND.n276 VGND.n275 0.141125
R6551 VGND.n91 VGND.n90 0.13201
R6552 VGND.n97 VGND.n96 0.13201
R6553 VGND.n103 VGND.n102 0.13201
R6554 VGND.n109 VGND.n108 0.13201
R6555 VGND.n115 VGND.n114 0.13201
R6556 VGND.n121 VGND.n120 0.13201
R6557 VGND.n127 VGND.n126 0.13201
R6558 VGND.n1772 VGND.n129 0.13201
R6559 VGND.n370 VGND.n341 0.13201
R6560 VGND.n374 VGND.n373 0.13201
R6561 VGND.n379 VGND.n378 0.13201
R6562 VGND.n385 VGND.n384 0.13201
R6563 VGND.n391 VGND.n390 0.13201
R6564 VGND.n397 VGND.n396 0.13201
R6565 VGND.n403 VGND.n402 0.13201
R6566 VGND.n409 VGND.n408 0.13201
R6567 VGND.n415 VGND.n414 0.13201
R6568 VGND.n421 VGND.n420 0.13201
R6569 VGND.n427 VGND.n426 0.13201
R6570 VGND.n433 VGND.n432 0.13201
R6571 VGND.n439 VGND.n438 0.13201
R6572 VGND.n445 VGND.n444 0.13201
R6573 VGND.n451 VGND.n450 0.13201
R6574 VGND.n457 VGND.n456 0.13201
R6575 VGND.n463 VGND.n462 0.13201
R6576 VGND.n469 VGND.n468 0.13201
R6577 VGND.n473 VGND.n472 0.13201
R6578 VGND.n23 VGND.n22 0.13201
R6579 VGND.n29 VGND.n28 0.13201
R6580 VGND.n35 VGND.n34 0.13201
R6581 VGND.n41 VGND.n40 0.13201
R6582 VGND.n47 VGND.n46 0.13201
R6583 VGND.n53 VGND.n52 0.13201
R6584 VGND.n59 VGND.n58 0.13201
R6585 VGND.n65 VGND.n64 0.13201
R6586 VGND.n1803 VGND.n67 0.13201
R6587 VGND.n741 VGND.n739 0.13201
R6588 VGND.n984 VGND.n983 0.13201
R6589 VGND.n964 VGND.n796 0.13201
R6590 VGND.n959 VGND.n799 0.13201
R6591 VGND.n942 VGND.n810 0.13201
R6592 VGND.n937 VGND.n813 0.13201
R6593 VGND.n920 VGND.n824 0.13201
R6594 VGND.n915 VGND.n827 0.13201
R6595 VGND.n898 VGND.n838 0.13201
R6596 VGND.n893 VGND.n841 0.13201
R6597 VGND.n876 VGND.n852 0.13201
R6598 VGND.n871 VGND.n855 0.13201
R6599 VGND.n148 VGND.n147 0.13201
R6600 VGND.n296 VGND.n295 0.13201
R6601 VGND.n290 VGND.n287 0.13201
R6602 VGND.n277 VGND.n276 0.13201
R6603 VGND.n271 VGND.n214 0.13201
R6604 VGND.n236 VGND.n0 0.13201
R6605 VGND.n996 VGND.n736 0.130708
R6606 VGND.n970 VGND.n969 0.130708
R6607 VGND.n947 VGND.n807 0.130708
R6608 VGND.n925 VGND.n821 0.130708
R6609 VGND.n903 VGND.n835 0.130708
R6610 VGND.n881 VGND.n849 0.130708
R6611 VGND.n181 VGND.n179 0.130708
R6612 VGND.n203 VGND.n202 0.130708
R6613 VGND.n594 VGND.n576 0.124275
R6614 VGND.n618 VGND.n598 0.124275
R6615 VGND.n642 VGND.n622 0.124275
R6616 VGND.n666 VGND.n646 0.124275
R6617 VGND.n690 VGND.n670 0.124275
R6618 VGND.n1064 VGND.n1063 0.124275
R6619 VGND.n1030 VGND.n707 0.124275
R6620 VGND.n1736 VGND.n1735 0.124275
R6621 VGND VGND.n1013 0.124198
R6622 VGND VGND.n981 0.124198
R6623 VGND VGND.n957 0.124198
R6624 VGND VGND.n935 0.124198
R6625 VGND VGND.n913 0.124198
R6626 VGND VGND.n891 0.124198
R6627 VGND VGND.n325 0.124198
R6628 VGND VGND.n198 0.124198
R6629 VGND.n1768 VGND.n1767 0.121824
R6630 VGND.n4 VGND.n2 0.121824
R6631 VGND.n1136 VGND.n1135 0.120598
R6632 VGND.n1123 VGND.n1122 0.120598
R6633 VGND.n1110 VGND.n1109 0.120598
R6634 VGND.n1097 VGND.n1096 0.120598
R6635 VGND.n1084 VGND.n1083 0.120598
R6636 VGND.n1065 VGND.n701 0.120598
R6637 VGND.n1058 VGND.n1057 0.120598
R6638 VGND.n1045 VGND.n338 0.120598
R6639 VGND.n1126 VGND 0.113245
R6640 VGND.n1113 VGND 0.113245
R6641 VGND.n1100 VGND 0.113245
R6642 VGND.n1087 VGND 0.113245
R6643 VGND.n1074 VGND 0.113245
R6644 VGND.n1061 VGND 0.113245
R6645 VGND.n1048 VGND 0.113245
R6646 VGND.n1733 VGND 0.113245
R6647 VGND.n1767 VGND.n1766 0.108343
R6648 VGND.n1834 VGND.n2 0.108343
R6649 VGND.n867 VGND.n866 0.104667
R6650 VGND.n863 VGND.n155 0.104667
R6651 VGND.n267 VGND.n219 0.104667
R6652 VGND.n248 VGND.n247 0.104667
R6653 VGND VGND.n1699 0.0721146
R6654 VGND.n1688 VGND 0.0721146
R6655 VGND VGND.n1681 0.0721146
R6656 VGND.n1670 VGND 0.0721146
R6657 VGND VGND.n1663 0.0721146
R6658 VGND VGND.n1644 0.0721146
R6659 VGND.n1772 VGND 0.0708125
R6660 VGND.n1803 VGND 0.0708125
R6661 VGND.n996 VGND 0.0695104
R6662 VGND.n969 VGND 0.0695104
R6663 VGND.n947 VGND 0.0695104
R6664 VGND.n925 VGND 0.0695104
R6665 VGND.n903 VGND 0.0695104
R6666 VGND.n881 VGND 0.0695104
R6667 VGND VGND.n181 0.0695104
R6668 VGND VGND.n203 0.0695104
R6669 VGND.n90 VGND.n87 0.0577917
R6670 VGND.n96 VGND.n92 0.0577917
R6671 VGND.n102 VGND.n98 0.0577917
R6672 VGND.n108 VGND.n104 0.0577917
R6673 VGND.n114 VGND.n110 0.0577917
R6674 VGND.n120 VGND.n116 0.0577917
R6675 VGND.n126 VGND.n122 0.0577917
R6676 VGND.n129 VGND.n128 0.0577917
R6677 VGND.n512 VGND.n341 0.0577917
R6678 VGND.n373 VGND.n372 0.0577917
R6679 VGND.n378 VGND.n375 0.0577917
R6680 VGND.n384 VGND.n380 0.0577917
R6681 VGND.n390 VGND.n386 0.0577917
R6682 VGND.n396 VGND.n392 0.0577917
R6683 VGND.n402 VGND.n398 0.0577917
R6684 VGND.n408 VGND.n404 0.0577917
R6685 VGND.n414 VGND.n410 0.0577917
R6686 VGND.n420 VGND.n416 0.0577917
R6687 VGND.n426 VGND.n422 0.0577917
R6688 VGND.n432 VGND.n428 0.0577917
R6689 VGND.n438 VGND.n434 0.0577917
R6690 VGND.n444 VGND.n440 0.0577917
R6691 VGND.n450 VGND.n446 0.0577917
R6692 VGND.n456 VGND.n452 0.0577917
R6693 VGND.n462 VGND.n458 0.0577917
R6694 VGND.n468 VGND.n464 0.0577917
R6695 VGND.n474 VGND.n473 0.0577917
R6696 VGND.n22 VGND.n19 0.0577917
R6697 VGND.n28 VGND.n24 0.0577917
R6698 VGND.n34 VGND.n30 0.0577917
R6699 VGND.n40 VGND.n36 0.0577917
R6700 VGND.n46 VGND.n42 0.0577917
R6701 VGND.n52 VGND.n48 0.0577917
R6702 VGND.n58 VGND.n54 0.0577917
R6703 VGND.n64 VGND.n60 0.0577917
R6704 VGND.n67 VGND.n66 0.0577917
R6705 VGND.n994 VGND.n739 0.0577917
R6706 VGND.n985 VGND.n984 0.0577917
R6707 VGND.n967 VGND.n796 0.0577917
R6708 VGND.n962 VGND.n799 0.0577917
R6709 VGND.n945 VGND.n810 0.0577917
R6710 VGND.n940 VGND.n813 0.0577917
R6711 VGND.n923 VGND.n824 0.0577917
R6712 VGND.n918 VGND.n827 0.0577917
R6713 VGND.n901 VGND.n838 0.0577917
R6714 VGND.n896 VGND.n841 0.0577917
R6715 VGND.n879 VGND.n852 0.0577917
R6716 VGND.n874 VGND.n855 0.0577917
R6717 VGND.n147 VGND.n143 0.0577917
R6718 VGND.n297 VGND.n296 0.0577917
R6719 VGND.n293 VGND.n287 0.0577917
R6720 VGND.n278 VGND.n277 0.0577917
R6721 VGND.n274 VGND.n214 0.0577917
R6722 VGND.n245 VGND.n236 0.0577917
R6723 VGND.n729 VGND 0.0522857
R6724 VGND.n172 VGND 0.0522857
R6725 VGND.n270 VGND 0.0213333
R6726 VGND VGND.n131 0.0164314
R6727 VGND VGND.n1835 0.0164314
R6728 VGND.n870 VGND 0.00918056
R6729 VGND.n270 VGND 0.00918056
R6730 VGND.n1014 VGND 0.00701042
R6731 VGND.n982 VGND 0.00701042
R6732 VGND.n958 VGND 0.00701042
R6733 VGND.n936 VGND 0.00701042
R6734 VGND.n914 VGND 0.00701042
R6735 VGND.n892 VGND 0.00701042
R6736 VGND.n326 VGND 0.00701042
R6737 VGND.n289 VGND 0.00701042
R6738 VGND.n1135 VGND.n576 0.00417647
R6739 VGND.n1122 VGND.n598 0.00417647
R6740 VGND.n1109 VGND.n622 0.00417647
R6741 VGND.n1096 VGND.n646 0.00417647
R6742 VGND.n1083 VGND.n670 0.00417647
R6743 VGND.n1065 VGND.n1064 0.00417647
R6744 VGND.n1057 VGND.n707 0.00417647
R6745 VGND.n1736 VGND.n338 0.00417647
R6746 a_9330_16954.n1 a_9330_16954.t9 543.053
R6747 a_9330_16954.n2 a_9330_16954.t29 543.053
R6748 a_9330_16954.n4 a_9330_16954.t16 543.053
R6749 a_9330_16954.n6 a_9330_16954.t35 543.053
R6750 a_9330_16954.n8 a_9330_16954.t23 543.053
R6751 a_9330_16954.n10 a_9330_16954.t25 543.053
R6752 a_9330_16954.n12 a_9330_16954.t11 543.053
R6753 a_9330_16954.n14 a_9330_16954.t31 543.053
R6754 a_9330_16954.n16 a_9330_16954.t19 543.053
R6755 a_9330_16954.n18 a_9330_16954.t37 543.053
R6756 a_9330_16954.n20 a_9330_16954.t18 543.053
R6757 a_9330_16954.n22 a_9330_16954.t36 543.053
R6758 a_9330_16954.n24 a_9330_16954.t24 543.053
R6759 a_9330_16954.n26 a_9330_16954.t10 543.053
R6760 a_9330_16954.n28 a_9330_16954.t30 543.053
R6761 a_9330_16954.n0 a_9330_16954.t17 543.053
R6762 a_9330_16954.n1 a_9330_16954.t38 221.72
R6763 a_9330_16954.n2 a_9330_16954.t26 221.72
R6764 a_9330_16954.n4 a_9330_16954.t12 221.72
R6765 a_9330_16954.n6 a_9330_16954.t32 221.72
R6766 a_9330_16954.n8 a_9330_16954.t20 221.72
R6767 a_9330_16954.n10 a_9330_16954.t22 221.72
R6768 a_9330_16954.n12 a_9330_16954.t8 221.72
R6769 a_9330_16954.n14 a_9330_16954.t28 221.72
R6770 a_9330_16954.n16 a_9330_16954.t15 221.72
R6771 a_9330_16954.n18 a_9330_16954.t34 221.72
R6772 a_9330_16954.n20 a_9330_16954.t14 221.72
R6773 a_9330_16954.n22 a_9330_16954.t33 221.72
R6774 a_9330_16954.n24 a_9330_16954.t21 221.72
R6775 a_9330_16954.n26 a_9330_16954.t39 221.72
R6776 a_9330_16954.n28 a_9330_16954.t27 221.72
R6777 a_9330_16954.n0 a_9330_16954.t13 221.72
R6778 a_9330_16954.n3 a_9330_16954.n1 218.32
R6779 a_9330_16954.n3 a_9330_16954.n2 217.734
R6780 a_9330_16954.n5 a_9330_16954.n4 217.734
R6781 a_9330_16954.n7 a_9330_16954.n6 217.734
R6782 a_9330_16954.n9 a_9330_16954.n8 217.734
R6783 a_9330_16954.n11 a_9330_16954.n10 217.734
R6784 a_9330_16954.n13 a_9330_16954.n12 217.734
R6785 a_9330_16954.n15 a_9330_16954.n14 217.734
R6786 a_9330_16954.n17 a_9330_16954.n16 217.734
R6787 a_9330_16954.n19 a_9330_16954.n18 217.734
R6788 a_9330_16954.n21 a_9330_16954.n20 217.734
R6789 a_9330_16954.n23 a_9330_16954.n22 217.734
R6790 a_9330_16954.n25 a_9330_16954.n24 217.734
R6791 a_9330_16954.n27 a_9330_16954.n26 217.734
R6792 a_9330_16954.n29 a_9330_16954.n28 217.734
R6793 a_9330_16954.n30 a_9330_16954.n0 213.234
R6794 a_9330_16954.n33 a_9330_16954.t6 85.2499
R6795 a_9330_16954.n35 a_9330_16954.t5 85.2499
R6796 a_9330_16954.t7 a_9330_16954.n37 85.2499
R6797 a_9330_16954.n31 a_9330_16954.t4 84.7173
R6798 a_9330_16954.n37 a_9330_16954.t3 83.7172
R6799 a_9330_16954.n32 a_9330_16954.t0 83.7172
R6800 a_9330_16954.n33 a_9330_16954.t2 83.7172
R6801 a_9330_16954.n35 a_9330_16954.t1 83.7172
R6802 a_9330_16954.n34 a_9330_16954.n32 5.16238
R6803 a_9330_16954.n36 a_9330_16954.n35 5.16238
R6804 a_9330_16954.n30 a_9330_16954.n29 5.08518
R6805 a_9330_16954.n34 a_9330_16954.n33 4.64452
R6806 a_9330_16954.n37 a_9330_16954.n36 4.64452
R6807 a_9330_16954.n5 a_9330_16954.n3 0.585177
R6808 a_9330_16954.n7 a_9330_16954.n5 0.585177
R6809 a_9330_16954.n9 a_9330_16954.n7 0.585177
R6810 a_9330_16954.n11 a_9330_16954.n9 0.585177
R6811 a_9330_16954.n13 a_9330_16954.n11 0.585177
R6812 a_9330_16954.n15 a_9330_16954.n13 0.585177
R6813 a_9330_16954.n17 a_9330_16954.n15 0.585177
R6814 a_9330_16954.n19 a_9330_16954.n17 0.585177
R6815 a_9330_16954.n21 a_9330_16954.n19 0.585177
R6816 a_9330_16954.n23 a_9330_16954.n21 0.585177
R6817 a_9330_16954.n25 a_9330_16954.n23 0.585177
R6818 a_9330_16954.n27 a_9330_16954.n25 0.585177
R6819 a_9330_16954.n29 a_9330_16954.n27 0.585177
R6820 a_9330_16954.n36 a_9330_16954.n34 0.518357
R6821 a_9330_16954.n32 a_9330_16954.n31 0.36463
R6822 a_9330_16954.n31 a_9330_16954.n30 0.226306
R6823 tdc_0.vernier_delay_line_0.stop_strong.n52 tdc_0.vernier_delay_line_0.stop_strong.t86 851.506
R6824 tdc_0.vernier_delay_line_0.stop_strong.n45 tdc_0.vernier_delay_line_0.stop_strong.t48 851.506
R6825 tdc_0.vernier_delay_line_0.stop_strong.n38 tdc_0.vernier_delay_line_0.stop_strong.t76 851.506
R6826 tdc_0.vernier_delay_line_0.stop_strong.n31 tdc_0.vernier_delay_line_0.stop_strong.t66 851.506
R6827 tdc_0.vernier_delay_line_0.stop_strong.n24 tdc_0.vernier_delay_line_0.stop_strong.t49 851.506
R6828 tdc_0.vernier_delay_line_0.stop_strong.n17 tdc_0.vernier_delay_line_0.stop_strong.t61 851.506
R6829 tdc_0.vernier_delay_line_0.stop_strong.n10 tdc_0.vernier_delay_line_0.stop_strong.t80 851.506
R6830 tdc_0.vernier_delay_line_0.stop_strong.n4 tdc_0.vernier_delay_line_0.stop_strong.t56 851.506
R6831 tdc_0.vernier_delay_line_0.stop_strong.n52 tdc_0.vernier_delay_line_0.stop_strong.t79 850.414
R6832 tdc_0.vernier_delay_line_0.stop_strong.n45 tdc_0.vernier_delay_line_0.stop_strong.t58 850.414
R6833 tdc_0.vernier_delay_line_0.stop_strong.n38 tdc_0.vernier_delay_line_0.stop_strong.t74 850.414
R6834 tdc_0.vernier_delay_line_0.stop_strong.n31 tdc_0.vernier_delay_line_0.stop_strong.t77 850.414
R6835 tdc_0.vernier_delay_line_0.stop_strong.n24 tdc_0.vernier_delay_line_0.stop_strong.t45 850.414
R6836 tdc_0.vernier_delay_line_0.stop_strong.n17 tdc_0.vernier_delay_line_0.stop_strong.t59 850.414
R6837 tdc_0.vernier_delay_line_0.stop_strong.n10 tdc_0.vernier_delay_line_0.stop_strong.t39 850.414
R6838 tdc_0.vernier_delay_line_0.stop_strong.n4 tdc_0.vernier_delay_line_0.stop_strong.t87 850.414
R6839 tdc_0.vernier_delay_line_0.stop_strong.n48 tdc_0.vernier_delay_line_0.stop_strong.t75 641.061
R6840 tdc_0.vernier_delay_line_0.stop_strong.n41 tdc_0.vernier_delay_line_0.stop_strong.t38 641.061
R6841 tdc_0.vernier_delay_line_0.stop_strong.n34 tdc_0.vernier_delay_line_0.stop_strong.t81 641.061
R6842 tdc_0.vernier_delay_line_0.stop_strong.n27 tdc_0.vernier_delay_line_0.stop_strong.t70 641.061
R6843 tdc_0.vernier_delay_line_0.stop_strong.n20 tdc_0.vernier_delay_line_0.stop_strong.t40 641.061
R6844 tdc_0.vernier_delay_line_0.stop_strong.n13 tdc_0.vernier_delay_line_0.stop_strong.t52 641.061
R6845 tdc_0.vernier_delay_line_0.stop_strong.n6 tdc_0.vernier_delay_line_0.stop_strong.t67 641.061
R6846 tdc_0.vernier_delay_line_0.stop_strong.n0 tdc_0.vernier_delay_line_0.stop_strong.t78 641.061
R6847 tdc_0.vernier_delay_line_0.stop_strong.n48 tdc_0.vernier_delay_line_0.stop_strong.t41 547.874
R6848 tdc_0.vernier_delay_line_0.stop_strong.n49 tdc_0.vernier_delay_line_0.stop_strong.t54 547.874
R6849 tdc_0.vernier_delay_line_0.stop_strong.n50 tdc_0.vernier_delay_line_0.stop_strong.t32 547.874
R6850 tdc_0.vernier_delay_line_0.stop_strong.n51 tdc_0.vernier_delay_line_0.stop_strong.t34 547.874
R6851 tdc_0.vernier_delay_line_0.stop_strong.n41 tdc_0.vernier_delay_line_0.stop_strong.t65 547.874
R6852 tdc_0.vernier_delay_line_0.stop_strong.n42 tdc_0.vernier_delay_line_0.stop_strong.t85 547.874
R6853 tdc_0.vernier_delay_line_0.stop_strong.n43 tdc_0.vernier_delay_line_0.stop_strong.t50 547.874
R6854 tdc_0.vernier_delay_line_0.stop_strong.n44 tdc_0.vernier_delay_line_0.stop_strong.t63 547.874
R6855 tdc_0.vernier_delay_line_0.stop_strong.n34 tdc_0.vernier_delay_line_0.stop_strong.t83 547.874
R6856 tdc_0.vernier_delay_line_0.stop_strong.n35 tdc_0.vernier_delay_line_0.stop_strong.t47 547.874
R6857 tdc_0.vernier_delay_line_0.stop_strong.n36 tdc_0.vernier_delay_line_0.stop_strong.t62 547.874
R6858 tdc_0.vernier_delay_line_0.stop_strong.n37 tdc_0.vernier_delay_line_0.stop_strong.t84 547.874
R6859 tdc_0.vernier_delay_line_0.stop_strong.n27 tdc_0.vernier_delay_line_0.stop_strong.t42 547.874
R6860 tdc_0.vernier_delay_line_0.stop_strong.n28 tdc_0.vernier_delay_line_0.stop_strong.t44 547.874
R6861 tdc_0.vernier_delay_line_0.stop_strong.n29 tdc_0.vernier_delay_line_0.stop_strong.t57 547.874
R6862 tdc_0.vernier_delay_line_0.stop_strong.n30 tdc_0.vernier_delay_line_0.stop_strong.t73 547.874
R6863 tdc_0.vernier_delay_line_0.stop_strong.n20 tdc_0.vernier_delay_line_0.stop_strong.t53 547.874
R6864 tdc_0.vernier_delay_line_0.stop_strong.n21 tdc_0.vernier_delay_line_0.stop_strong.t69 547.874
R6865 tdc_0.vernier_delay_line_0.stop_strong.n22 tdc_0.vernier_delay_line_0.stop_strong.t71 547.874
R6866 tdc_0.vernier_delay_line_0.stop_strong.n23 tdc_0.vernier_delay_line_0.stop_strong.t36 547.874
R6867 tdc_0.vernier_delay_line_0.stop_strong.n13 tdc_0.vernier_delay_line_0.stop_strong.t68 547.874
R6868 tdc_0.vernier_delay_line_0.stop_strong.n14 tdc_0.vernier_delay_line_0.stop_strong.t35 547.874
R6869 tdc_0.vernier_delay_line_0.stop_strong.n15 tdc_0.vernier_delay_line_0.stop_strong.t51 547.874
R6870 tdc_0.vernier_delay_line_0.stop_strong.n16 tdc_0.vernier_delay_line_0.stop_strong.t64 547.874
R6871 tdc_0.vernier_delay_line_0.stop_strong.n6 tdc_0.vernier_delay_line_0.stop_strong.t33 547.874
R6872 tdc_0.vernier_delay_line_0.stop_strong.n7 tdc_0.vernier_delay_line_0.stop_strong.t60 547.874
R6873 tdc_0.vernier_delay_line_0.stop_strong.n8 tdc_0.vernier_delay_line_0.stop_strong.t82 547.874
R6874 tdc_0.vernier_delay_line_0.stop_strong.n9 tdc_0.vernier_delay_line_0.stop_strong.t46 547.874
R6875 tdc_0.vernier_delay_line_0.stop_strong.n0 tdc_0.vernier_delay_line_0.stop_strong.t43 547.874
R6876 tdc_0.vernier_delay_line_0.stop_strong.n1 tdc_0.vernier_delay_line_0.stop_strong.t55 547.874
R6877 tdc_0.vernier_delay_line_0.stop_strong.n2 tdc_0.vernier_delay_line_0.stop_strong.t72 547.874
R6878 tdc_0.vernier_delay_line_0.stop_strong.n3 tdc_0.vernier_delay_line_0.stop_strong.t37 547.874
R6879 tdc_0.vernier_delay_line_0.stop_strong.n53 tdc_0.vernier_delay_line_0.stop_strong.n51 189.41
R6880 tdc_0.vernier_delay_line_0.stop_strong.n46 tdc_0.vernier_delay_line_0.stop_strong.n44 189.41
R6881 tdc_0.vernier_delay_line_0.stop_strong.n39 tdc_0.vernier_delay_line_0.stop_strong.n37 189.41
R6882 tdc_0.vernier_delay_line_0.stop_strong.n32 tdc_0.vernier_delay_line_0.stop_strong.n30 189.41
R6883 tdc_0.vernier_delay_line_0.stop_strong.n25 tdc_0.vernier_delay_line_0.stop_strong.n23 189.41
R6884 tdc_0.vernier_delay_line_0.stop_strong.n18 tdc_0.vernier_delay_line_0.stop_strong.n16 189.41
R6885 tdc_0.vernier_delay_line_0.stop_strong.n11 tdc_0.vernier_delay_line_0.stop_strong.n9 189.41
R6886 tdc_0.vernier_delay_line_0.stop_strong.n5 tdc_0.vernier_delay_line_0.stop_strong.n3 189.41
R6887 tdc_0.vernier_delay_line_0.stop_strong.n49 tdc_0.vernier_delay_line_0.stop_strong.n48 93.1872
R6888 tdc_0.vernier_delay_line_0.stop_strong.n50 tdc_0.vernier_delay_line_0.stop_strong.n49 93.1872
R6889 tdc_0.vernier_delay_line_0.stop_strong.n51 tdc_0.vernier_delay_line_0.stop_strong.n50 93.1872
R6890 tdc_0.vernier_delay_line_0.stop_strong.n42 tdc_0.vernier_delay_line_0.stop_strong.n41 93.1872
R6891 tdc_0.vernier_delay_line_0.stop_strong.n43 tdc_0.vernier_delay_line_0.stop_strong.n42 93.1872
R6892 tdc_0.vernier_delay_line_0.stop_strong.n44 tdc_0.vernier_delay_line_0.stop_strong.n43 93.1872
R6893 tdc_0.vernier_delay_line_0.stop_strong.n35 tdc_0.vernier_delay_line_0.stop_strong.n34 93.1872
R6894 tdc_0.vernier_delay_line_0.stop_strong.n36 tdc_0.vernier_delay_line_0.stop_strong.n35 93.1872
R6895 tdc_0.vernier_delay_line_0.stop_strong.n37 tdc_0.vernier_delay_line_0.stop_strong.n36 93.1872
R6896 tdc_0.vernier_delay_line_0.stop_strong.n28 tdc_0.vernier_delay_line_0.stop_strong.n27 93.1872
R6897 tdc_0.vernier_delay_line_0.stop_strong.n29 tdc_0.vernier_delay_line_0.stop_strong.n28 93.1872
R6898 tdc_0.vernier_delay_line_0.stop_strong.n30 tdc_0.vernier_delay_line_0.stop_strong.n29 93.1872
R6899 tdc_0.vernier_delay_line_0.stop_strong.n21 tdc_0.vernier_delay_line_0.stop_strong.n20 93.1872
R6900 tdc_0.vernier_delay_line_0.stop_strong.n22 tdc_0.vernier_delay_line_0.stop_strong.n21 93.1872
R6901 tdc_0.vernier_delay_line_0.stop_strong.n23 tdc_0.vernier_delay_line_0.stop_strong.n22 93.1872
R6902 tdc_0.vernier_delay_line_0.stop_strong.n14 tdc_0.vernier_delay_line_0.stop_strong.n13 93.1872
R6903 tdc_0.vernier_delay_line_0.stop_strong.n15 tdc_0.vernier_delay_line_0.stop_strong.n14 93.1872
R6904 tdc_0.vernier_delay_line_0.stop_strong.n16 tdc_0.vernier_delay_line_0.stop_strong.n15 93.1872
R6905 tdc_0.vernier_delay_line_0.stop_strong.n7 tdc_0.vernier_delay_line_0.stop_strong.n6 93.1872
R6906 tdc_0.vernier_delay_line_0.stop_strong.n8 tdc_0.vernier_delay_line_0.stop_strong.n7 93.1872
R6907 tdc_0.vernier_delay_line_0.stop_strong.n9 tdc_0.vernier_delay_line_0.stop_strong.n8 93.1872
R6908 tdc_0.vernier_delay_line_0.stop_strong.n1 tdc_0.vernier_delay_line_0.stop_strong.n0 93.1872
R6909 tdc_0.vernier_delay_line_0.stop_strong.n2 tdc_0.vernier_delay_line_0.stop_strong.n1 93.1872
R6910 tdc_0.vernier_delay_line_0.stop_strong.n3 tdc_0.vernier_delay_line_0.stop_strong.n2 93.1872
R6911 tdc_0.vernier_delay_line_0.stop_strong.n82 tdc_0.vernier_delay_line_0.stop_strong.t21 85.2499
R6912 tdc_0.vernier_delay_line_0.stop_strong.n80 tdc_0.vernier_delay_line_0.stop_strong.t28 85.2499
R6913 tdc_0.vernier_delay_line_0.stop_strong.n78 tdc_0.vernier_delay_line_0.stop_strong.t18 85.2499
R6914 tdc_0.vernier_delay_line_0.stop_strong.n76 tdc_0.vernier_delay_line_0.stop_strong.t24 85.2499
R6915 tdc_0.vernier_delay_line_0.stop_strong.n74 tdc_0.vernier_delay_line_0.stop_strong.t22 85.2499
R6916 tdc_0.vernier_delay_line_0.stop_strong.n72 tdc_0.vernier_delay_line_0.stop_strong.t29 85.2499
R6917 tdc_0.vernier_delay_line_0.stop_strong.n70 tdc_0.vernier_delay_line_0.stop_strong.t19 85.2499
R6918 tdc_0.vernier_delay_line_0.stop_strong.n68 tdc_0.vernier_delay_line_0.stop_strong.t25 85.2499
R6919 tdc_0.vernier_delay_line_0.stop_strong.n66 tdc_0.vernier_delay_line_0.stop_strong.t16 85.2499
R6920 tdc_0.vernier_delay_line_0.stop_strong.n64 tdc_0.vernier_delay_line_0.stop_strong.t26 85.2499
R6921 tdc_0.vernier_delay_line_0.stop_strong.n62 tdc_0.vernier_delay_line_0.stop_strong.t17 85.2499
R6922 tdc_0.vernier_delay_line_0.stop_strong.n60 tdc_0.vernier_delay_line_0.stop_strong.t23 85.2499
R6923 tdc_0.vernier_delay_line_0.stop_strong.n58 tdc_0.vernier_delay_line_0.stop_strong.t30 85.2499
R6924 tdc_0.vernier_delay_line_0.stop_strong.n56 tdc_0.vernier_delay_line_0.stop_strong.t20 85.2499
R6925 tdc_0.vernier_delay_line_0.stop_strong.n55 tdc_0.vernier_delay_line_0.stop_strong.t27 85.2499
R6926 tdc_0.vernier_delay_line_0.stop_strong.n86 tdc_0.vernier_delay_line_0.stop_strong.t31 84.7281
R6927 tdc_0.vernier_delay_line_0.stop_strong.n85 tdc_0.vernier_delay_line_0.stop_strong.t1 83.7172
R6928 tdc_0.vernier_delay_line_0.stop_strong.n82 tdc_0.vernier_delay_line_0.stop_strong.t7 83.7172
R6929 tdc_0.vernier_delay_line_0.stop_strong.n80 tdc_0.vernier_delay_line_0.stop_strong.t14 83.7172
R6930 tdc_0.vernier_delay_line_0.stop_strong.n78 tdc_0.vernier_delay_line_0.stop_strong.t4 83.7172
R6931 tdc_0.vernier_delay_line_0.stop_strong.n76 tdc_0.vernier_delay_line_0.stop_strong.t10 83.7172
R6932 tdc_0.vernier_delay_line_0.stop_strong.n74 tdc_0.vernier_delay_line_0.stop_strong.t8 83.7172
R6933 tdc_0.vernier_delay_line_0.stop_strong.n72 tdc_0.vernier_delay_line_0.stop_strong.t15 83.7172
R6934 tdc_0.vernier_delay_line_0.stop_strong.n70 tdc_0.vernier_delay_line_0.stop_strong.t5 83.7172
R6935 tdc_0.vernier_delay_line_0.stop_strong.n68 tdc_0.vernier_delay_line_0.stop_strong.t11 83.7172
R6936 tdc_0.vernier_delay_line_0.stop_strong.n66 tdc_0.vernier_delay_line_0.stop_strong.t2 83.7172
R6937 tdc_0.vernier_delay_line_0.stop_strong.n64 tdc_0.vernier_delay_line_0.stop_strong.t12 83.7172
R6938 tdc_0.vernier_delay_line_0.stop_strong.n62 tdc_0.vernier_delay_line_0.stop_strong.t3 83.7172
R6939 tdc_0.vernier_delay_line_0.stop_strong.n60 tdc_0.vernier_delay_line_0.stop_strong.t9 83.7172
R6940 tdc_0.vernier_delay_line_0.stop_strong.n58 tdc_0.vernier_delay_line_0.stop_strong.t0 83.7172
R6941 tdc_0.vernier_delay_line_0.stop_strong.n56 tdc_0.vernier_delay_line_0.stop_strong.t6 83.7172
R6942 tdc_0.vernier_delay_line_0.stop_strong.n55 tdc_0.vernier_delay_line_0.stop_strong.t13 83.7172
R6943 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n5 11.8482
R6944 tdc_0.vernier_delay_line_0.stop_strong.n54 tdc_0.vernier_delay_line_0.stop_strong.n53 9.66066
R6945 tdc_0.vernier_delay_line_0.stop_strong.n47 tdc_0.vernier_delay_line_0.stop_strong.n46 9.66066
R6946 tdc_0.vernier_delay_line_0.stop_strong.n40 tdc_0.vernier_delay_line_0.stop_strong.n39 9.66066
R6947 tdc_0.vernier_delay_line_0.stop_strong.n33 tdc_0.vernier_delay_line_0.stop_strong.n32 9.66066
R6948 tdc_0.vernier_delay_line_0.stop_strong.n26 tdc_0.vernier_delay_line_0.stop_strong.n25 9.66066
R6949 tdc_0.vernier_delay_line_0.stop_strong.n19 tdc_0.vernier_delay_line_0.stop_strong.n18 9.66066
R6950 tdc_0.vernier_delay_line_0.stop_strong.n12 tdc_0.vernier_delay_line_0.stop_strong.n11 9.66066
R6951 tdc_0.vernier_delay_line_0.stop_strong.n84 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk 8.04701
R6952 tdc_0.vernier_delay_line_0.stop_strong.n57 tdc_0.vernier_delay_line_0.stop_strong.n55 5.16238
R6953 tdc_0.vernier_delay_line_0.stop_strong.n83 tdc_0.vernier_delay_line_0.stop_strong.n82 4.64452
R6954 tdc_0.vernier_delay_line_0.stop_strong.n81 tdc_0.vernier_delay_line_0.stop_strong.n80 4.64452
R6955 tdc_0.vernier_delay_line_0.stop_strong.n79 tdc_0.vernier_delay_line_0.stop_strong.n78 4.64452
R6956 tdc_0.vernier_delay_line_0.stop_strong.n77 tdc_0.vernier_delay_line_0.stop_strong.n76 4.64452
R6957 tdc_0.vernier_delay_line_0.stop_strong.n75 tdc_0.vernier_delay_line_0.stop_strong.n74 4.64452
R6958 tdc_0.vernier_delay_line_0.stop_strong.n73 tdc_0.vernier_delay_line_0.stop_strong.n72 4.64452
R6959 tdc_0.vernier_delay_line_0.stop_strong.n71 tdc_0.vernier_delay_line_0.stop_strong.n70 4.64452
R6960 tdc_0.vernier_delay_line_0.stop_strong.n69 tdc_0.vernier_delay_line_0.stop_strong.n68 4.64452
R6961 tdc_0.vernier_delay_line_0.stop_strong.n67 tdc_0.vernier_delay_line_0.stop_strong.n66 4.64452
R6962 tdc_0.vernier_delay_line_0.stop_strong.n65 tdc_0.vernier_delay_line_0.stop_strong.n64 4.64452
R6963 tdc_0.vernier_delay_line_0.stop_strong.n63 tdc_0.vernier_delay_line_0.stop_strong.n62 4.64452
R6964 tdc_0.vernier_delay_line_0.stop_strong.n61 tdc_0.vernier_delay_line_0.stop_strong.n60 4.64452
R6965 tdc_0.vernier_delay_line_0.stop_strong.n59 tdc_0.vernier_delay_line_0.stop_strong.n58 4.64452
R6966 tdc_0.vernier_delay_line_0.stop_strong.n57 tdc_0.vernier_delay_line_0.stop_strong.n56 4.64452
R6967 tdc_0.vernier_delay_line_0.stop_strong.n85 tdc_0.vernier_delay_line_0.stop_strong.n84 4.64452
R6968 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n12 2.188
R6969 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n19 2.188
R6970 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n26 2.188
R6971 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n33 2.188
R6972 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n40 2.188
R6973 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n47 2.188
R6974 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk tdc_0.vernier_delay_line_0.stop_strong.n54 2.188
R6975 tdc_0.vernier_delay_line_0.stop_strong.n53 tdc_0.vernier_delay_line_0.stop_strong.n52 1.05649
R6976 tdc_0.vernier_delay_line_0.stop_strong.n46 tdc_0.vernier_delay_line_0.stop_strong.n45 1.05649
R6977 tdc_0.vernier_delay_line_0.stop_strong.n39 tdc_0.vernier_delay_line_0.stop_strong.n38 1.05649
R6978 tdc_0.vernier_delay_line_0.stop_strong.n32 tdc_0.vernier_delay_line_0.stop_strong.n31 1.05649
R6979 tdc_0.vernier_delay_line_0.stop_strong.n25 tdc_0.vernier_delay_line_0.stop_strong.n24 1.05649
R6980 tdc_0.vernier_delay_line_0.stop_strong.n18 tdc_0.vernier_delay_line_0.stop_strong.n17 1.05649
R6981 tdc_0.vernier_delay_line_0.stop_strong.n11 tdc_0.vernier_delay_line_0.stop_strong.n10 1.05649
R6982 tdc_0.vernier_delay_line_0.stop_strong.n5 tdc_0.vernier_delay_line_0.stop_strong.n4 1.05649
R6983 tdc_0.vernier_delay_line_0.stop_strong.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk 0.6655
R6984 tdc_0.vernier_delay_line_0.stop_strong.n19 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk 0.6655
R6985 tdc_0.vernier_delay_line_0.stop_strong.n26 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk 0.6655
R6986 tdc_0.vernier_delay_line_0.stop_strong.n33 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk 0.6655
R6987 tdc_0.vernier_delay_line_0.stop_strong.n40 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk 0.6655
R6988 tdc_0.vernier_delay_line_0.stop_strong.n47 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk 0.6655
R6989 tdc_0.vernier_delay_line_0.stop_strong.n54 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk 0.6655
R6990 tdc_0.vernier_delay_line_0.stop_strong.n83 tdc_0.vernier_delay_line_0.stop_strong.n81 0.518357
R6991 tdc_0.vernier_delay_line_0.stop_strong.n81 tdc_0.vernier_delay_line_0.stop_strong.n79 0.518357
R6992 tdc_0.vernier_delay_line_0.stop_strong.n79 tdc_0.vernier_delay_line_0.stop_strong.n77 0.518357
R6993 tdc_0.vernier_delay_line_0.stop_strong.n77 tdc_0.vernier_delay_line_0.stop_strong.n75 0.518357
R6994 tdc_0.vernier_delay_line_0.stop_strong.n75 tdc_0.vernier_delay_line_0.stop_strong.n73 0.518357
R6995 tdc_0.vernier_delay_line_0.stop_strong.n73 tdc_0.vernier_delay_line_0.stop_strong.n71 0.518357
R6996 tdc_0.vernier_delay_line_0.stop_strong.n71 tdc_0.vernier_delay_line_0.stop_strong.n69 0.518357
R6997 tdc_0.vernier_delay_line_0.stop_strong.n69 tdc_0.vernier_delay_line_0.stop_strong.n67 0.518357
R6998 tdc_0.vernier_delay_line_0.stop_strong.n67 tdc_0.vernier_delay_line_0.stop_strong.n65 0.518357
R6999 tdc_0.vernier_delay_line_0.stop_strong.n65 tdc_0.vernier_delay_line_0.stop_strong.n63 0.518357
R7000 tdc_0.vernier_delay_line_0.stop_strong.n63 tdc_0.vernier_delay_line_0.stop_strong.n61 0.518357
R7001 tdc_0.vernier_delay_line_0.stop_strong.n61 tdc_0.vernier_delay_line_0.stop_strong.n59 0.518357
R7002 tdc_0.vernier_delay_line_0.stop_strong.n59 tdc_0.vernier_delay_line_0.stop_strong.n57 0.518357
R7003 tdc_0.vernier_delay_line_0.stop_strong.n84 tdc_0.vernier_delay_line_0.stop_strong.n83 0.497131
R7004 tdc_0.vernier_delay_line_0.stop_strong.n86 tdc_0.vernier_delay_line_0.stop_strong.n85 0.3755
R7005 tdc_0.stop_buffer_0.stop_strong tdc_0.vernier_delay_line_0.stop_strong.n86 0.234296
R7006 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 784.053
R7007 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 784.053
R7008 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 784.053
R7009 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 784.053
R7010 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 539.841
R7011 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 539.841
R7012 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 539.841
R7013 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 539.841
R7014 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 215.293
R7015 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 215.293
R7016 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 215.293
R7017 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 215.293
R7018 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 168.659
R7019 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 167.992
R7020 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 166.144
R7021 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 165.8
R7022 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 85.2499
R7023 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 85.2499
R7024 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 83.7172
R7025 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 83.7172
R7026 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 75.7282
R7027 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 66.3172
R7028 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 36.1505
R7029 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 36.1505
R7030 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 34.5438
R7031 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 34.5438
R7032 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 17.4005
R7033 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 17.4005
R7034 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 17.2391
R7035 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 9.52217
R7036 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 9.52217
R7037 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 6.39571
R7038 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 5.30824
R7039 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 4.94887
R7040 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd 1.64112
R7041 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 1.06691
R7042 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 0.930188
R7043 a_10108_39954.n2 a_10108_39954.n1 34.9195
R7044 a_10108_39954.n3 a_10108_39954.n2 25.5407
R7045 a_10108_39954.n2 a_10108_39954.n0 25.2907
R7046 a_10108_39954.n1 a_10108_39954.t4 5.8005
R7047 a_10108_39954.n1 a_10108_39954.t5 5.8005
R7048 a_10108_39954.n0 a_10108_39954.t3 5.8005
R7049 a_10108_39954.n0 a_10108_39954.t2 5.8005
R7050 a_10108_39954.t0 a_10108_39954.n3 5.8005
R7051 a_10108_39954.n3 a_10108_39954.t1 5.8005
R7052 a_10958_39338.n1 a_10958_39338.t1 31.9657
R7053 a_10958_39338.n1 a_10958_39338.n0 25.8125
R7054 a_10958_39338.n3 a_10958_39338.n2 25.8125
R7055 a_10958_39338.n5 a_10958_39338.n4 25.8125
R7056 a_10958_39338.n10 a_10958_39338.n9 25.7038
R7057 a_10958_39338.n9 a_10958_39338.n8 25.3505
R7058 a_10958_39338.n7 a_10958_39338.n6 24.288
R7059 a_10958_39338.n6 a_10958_39338.t2 5.8005
R7060 a_10958_39338.n6 a_10958_39338.t10 5.8005
R7061 a_10958_39338.n0 a_10958_39338.t8 5.8005
R7062 a_10958_39338.n0 a_10958_39338.t0 5.8005
R7063 a_10958_39338.n2 a_10958_39338.t12 5.8005
R7064 a_10958_39338.n2 a_10958_39338.t11 5.8005
R7065 a_10958_39338.n4 a_10958_39338.t9 5.8005
R7066 a_10958_39338.n4 a_10958_39338.t7 5.8005
R7067 a_10958_39338.n8 a_10958_39338.t4 5.8005
R7068 a_10958_39338.n8 a_10958_39338.t5 5.8005
R7069 a_10958_39338.t6 a_10958_39338.n10 5.8005
R7070 a_10958_39338.n10 a_10958_39338.t3 5.8005
R7071 a_10958_39338.n7 a_10958_39338.n5 1.87822
R7072 a_10958_39338.n9 a_10958_39338.n7 1.41626
R7073 a_10958_39338.n3 a_10958_39338.n1 0.353761
R7074 a_10958_39338.n5 a_10958_39338.n3 0.353761
R7075 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 890.727
R7076 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 742.783
R7077 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 641.061
R7078 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 623.388
R7079 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 547.874
R7080 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 431.807
R7081 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 427.875
R7082 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7083 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7084 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7085 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7086 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 31.2103
R7087 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 31.0962
R7088 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 9.52217
R7089 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R7090 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 8.91506
R7091 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7092 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7093 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7094 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7095 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 879.481
R7096 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 742.783
R7097 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 641.061
R7098 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 623.388
R7099 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 547.874
R7100 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 431.807
R7101 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 427.875
R7102 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 333.161
R7103 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7104 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 168.077
R7105 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 75.5951
R7106 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R7107 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 31.2972
R7108 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 11.1806
R7109 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7110 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7111 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R7112 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7113 a_10108_28544.n2 a_10108_28544.n1 34.9195
R7114 a_10108_28544.n3 a_10108_28544.n2 25.5407
R7115 a_10108_28544.n2 a_10108_28544.n0 25.2907
R7116 a_10108_28544.n1 a_10108_28544.t4 5.8005
R7117 a_10108_28544.n1 a_10108_28544.t2 5.8005
R7118 a_10108_28544.n0 a_10108_28544.t3 5.8005
R7119 a_10108_28544.n0 a_10108_28544.t5 5.8005
R7120 a_10108_28544.n3 a_10108_28544.t0 5.8005
R7121 a_10108_28544.t1 a_10108_28544.n3 5.8005
R7122 a_10958_23364.n1 a_10958_23364.t1 31.9657
R7123 a_10958_23364.n1 a_10958_23364.n0 25.8125
R7124 a_10958_23364.n3 a_10958_23364.n2 25.8125
R7125 a_10958_23364.n5 a_10958_23364.n4 25.8125
R7126 a_10958_23364.n10 a_10958_23364.n9 25.7038
R7127 a_10958_23364.n9 a_10958_23364.n8 25.3505
R7128 a_10958_23364.n7 a_10958_23364.n6 24.288
R7129 a_10958_23364.n6 a_10958_23364.t2 5.8005
R7130 a_10958_23364.n6 a_10958_23364.t7 5.8005
R7131 a_10958_23364.n0 a_10958_23364.t10 5.8005
R7132 a_10958_23364.n0 a_10958_23364.t11 5.8005
R7133 a_10958_23364.n2 a_10958_23364.t12 5.8005
R7134 a_10958_23364.n2 a_10958_23364.t9 5.8005
R7135 a_10958_23364.n4 a_10958_23364.t8 5.8005
R7136 a_10958_23364.n4 a_10958_23364.t0 5.8005
R7137 a_10958_23364.n8 a_10958_23364.t3 5.8005
R7138 a_10958_23364.n8 a_10958_23364.t4 5.8005
R7139 a_10958_23364.n10 a_10958_23364.t5 5.8005
R7140 a_10958_23364.t6 a_10958_23364.n10 5.8005
R7141 a_10958_23364.n7 a_10958_23364.n5 1.87822
R7142 a_10958_23364.n9 a_10958_23364.n7 1.41626
R7143 a_10958_23364.n3 a_10958_23364.n1 0.353761
R7144 a_10958_23364.n5 a_10958_23364.n3 0.353761
R7145 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t2 628.097
R7146 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t6 622.766
R7147 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t4 523.774
R7148 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t5 304.647
R7149 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t7 304.647
R7150 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t3 202.44
R7151 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 169.062
R7152 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 166.237
R7153 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t0 84.7557
R7154 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t1 84.1197
R7155 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 12.6535
R7156 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 5.48979
R7157 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 4.5005
R7158 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 1.09595
R7159 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 879.481
R7160 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 742.783
R7161 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 641.061
R7162 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 623.388
R7163 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 547.874
R7164 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 431.807
R7165 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 427.875
R7166 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 333.161
R7167 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7168 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 168.077
R7169 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 75.5951
R7170 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 31.2972
R7171 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R7172 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 11.1806
R7173 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7174 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R7175 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7176 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7177 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 890.727
R7178 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 742.783
R7179 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 641.061
R7180 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 623.388
R7181 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 547.874
R7182 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 431.807
R7183 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 427.875
R7184 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7185 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7186 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7187 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7188 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 31.2103
R7189 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 31.0962
R7190 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R7191 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7192 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 8.91506
R7193 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7194 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7195 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7196 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7197 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 879.481
R7198 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 742.783
R7199 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 641.061
R7200 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 623.388
R7201 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 547.874
R7202 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 431.807
R7203 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 427.875
R7204 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 333.161
R7205 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7206 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 168.077
R7207 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 75.5951
R7208 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R7209 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R7210 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 11.1806
R7211 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7212 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7213 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R7214 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7215 a_10108_35390.n2 a_10108_35390.n1 34.9195
R7216 a_10108_35390.n3 a_10108_35390.n2 25.5407
R7217 a_10108_35390.n2 a_10108_35390.n0 25.2907
R7218 a_10108_35390.n1 a_10108_35390.t2 5.8005
R7219 a_10108_35390.n1 a_10108_35390.t5 5.8005
R7220 a_10108_35390.n0 a_10108_35390.t4 5.8005
R7221 a_10108_35390.n0 a_10108_35390.t3 5.8005
R7222 a_10108_35390.n3 a_10108_35390.t0 5.8005
R7223 a_10108_35390.t1 a_10108_35390.n3 5.8005
R7224 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 879.481
R7225 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 742.783
R7226 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 641.061
R7227 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 623.388
R7228 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 547.874
R7229 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 431.807
R7230 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 427.875
R7231 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 333.161
R7232 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7233 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 168.077
R7234 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 75.5951
R7235 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 31.2972
R7236 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R7237 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 11.1806
R7238 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7239 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7240 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R7241 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7242 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 890.727
R7243 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 742.783
R7244 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 641.061
R7245 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 623.388
R7246 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 547.874
R7247 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 431.807
R7248 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 427.875
R7249 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7250 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7251 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7252 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7253 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 31.2103
R7254 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 31.0962
R7255 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7256 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R7257 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 8.91506
R7258 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7259 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7260 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7261 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7262 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t4 628.097
R7263 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t7 622.766
R7264 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t5 523.774
R7265 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t6 304.647
R7266 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t2 304.647
R7267 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t3 202.44
R7268 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 169.062
R7269 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 166.237
R7270 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t0 84.7557
R7271 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t1 84.1197
R7272 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 12.6535
R7273 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 5.48979
R7274 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 4.5005
R7275 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 1.09595
R7276 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 552.84
R7277 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 552.84
R7278 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 552.84
R7279 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 552.84
R7280 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 539.841
R7281 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 539.841
R7282 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 539.841
R7283 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 539.841
R7284 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 215.293
R7285 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 215.293
R7286 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 215.293
R7287 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 215.293
R7288 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 166.468
R7289 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 166.149
R7290 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 165.8
R7291 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 165.8
R7292 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 85.1574
R7293 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 83.8097
R7294 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 83.8097
R7295 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 83.7172
R7296 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 74.288
R7297 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 67.7574
R7298 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 36.1505
R7299 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 36.1505
R7300 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 34.5438
R7301 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 34.5438
R7302 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 17.4005
R7303 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 17.4005
R7304 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 16.09
R7305 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 11.8364
R7306 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 9.52217
R7307 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 9.52217
R7308 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d 5.96628
R7309 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 5.83219
R7310 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 5.74235
R7311 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 5.49235
R7312 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 2.48878
R7313 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 1.44072
R7314 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 1.32081
R7315 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t6 628.097
R7316 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t4 622.766
R7317 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t2 523.774
R7318 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t3 304.647
R7319 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t5 304.647
R7320 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t7 202.44
R7321 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 169.062
R7322 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 166.237
R7323 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t1 84.7557
R7324 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t0 84.1197
R7325 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 12.6535
R7326 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 5.48979
R7327 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 4.5005
R7328 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 1.09595
R7329 a_10958_37056.n2 a_10958_37056.t4 31.9657
R7330 a_10958_37056.n2 a_10958_37056.n1 25.8125
R7331 a_10958_37056.n4 a_10958_37056.n3 25.8125
R7332 a_10958_37056.n6 a_10958_37056.n5 25.8125
R7333 a_10958_37056.n9 a_10958_37056.n0 25.7038
R7334 a_10958_37056.n10 a_10958_37056.n9 25.3505
R7335 a_10958_37056.n8 a_10958_37056.n7 24.288
R7336 a_10958_37056.n7 a_10958_37056.t7 5.8005
R7337 a_10958_37056.n7 a_10958_37056.t0 5.8005
R7338 a_10958_37056.n1 a_10958_37056.t2 5.8005
R7339 a_10958_37056.n1 a_10958_37056.t12 5.8005
R7340 a_10958_37056.n3 a_10958_37056.t5 5.8005
R7341 a_10958_37056.n3 a_10958_37056.t3 5.8005
R7342 a_10958_37056.n5 a_10958_37056.t11 5.8005
R7343 a_10958_37056.n5 a_10958_37056.t1 5.8005
R7344 a_10958_37056.n0 a_10958_37056.t9 5.8005
R7345 a_10958_37056.n0 a_10958_37056.t6 5.8005
R7346 a_10958_37056.n10 a_10958_37056.t8 5.8005
R7347 a_10958_37056.t10 a_10958_37056.n10 5.8005
R7348 a_10958_37056.n8 a_10958_37056.n6 1.87822
R7349 a_10958_37056.n9 a_10958_37056.n8 1.41626
R7350 a_10958_37056.n4 a_10958_37056.n2 0.353761
R7351 a_10958_37056.n6 a_10958_37056.n4 0.353761
R7352 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 890.727
R7353 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 742.783
R7354 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 641.061
R7355 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 623.388
R7356 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 547.874
R7357 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 431.807
R7358 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 427.875
R7359 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7360 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7361 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7362 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7363 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 31.2103
R7364 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 31.0962
R7365 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R7366 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7367 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 8.91506
R7368 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7369 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7370 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7371 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7372 a_10108_26262.n2 a_10108_26262.n1 34.9195
R7373 a_10108_26262.n3 a_10108_26262.n2 25.5407
R7374 a_10108_26262.n2 a_10108_26262.n0 25.2907
R7375 a_10108_26262.n1 a_10108_26262.t1 5.8005
R7376 a_10108_26262.n1 a_10108_26262.t0 5.8005
R7377 a_10108_26262.n0 a_10108_26262.t3 5.8005
R7378 a_10108_26262.n0 a_10108_26262.t2 5.8005
R7379 a_10108_26262.n3 a_10108_26262.t5 5.8005
R7380 a_10108_26262.t4 a_10108_26262.n3 5.8005
R7381 uo_out[6].n0 uo_out[6].t5 734.539
R7382 uo_out[6].n0 uo_out[6].t4 233.26
R7383 uo_out[6].n2 uo_out[6].n0 162.335
R7384 uo_out[6].n2 uo_out[6].n1 75.5733
R7385 uo_out[6].n4 uo_out[6].n3 66.3172
R7386 uo_out[6].n3 uo_out[6].t1 17.4005
R7387 uo_out[6].n3 uo_out[6].t3 17.4005
R7388 uo_out[6].n5 uo_out[6] 16.4025
R7389 uo_out[6].n1 uo_out[6].t2 9.52217
R7390 uo_out[6].n1 uo_out[6].t0 9.52217
R7391 uo_out[6].n5 uo_out[6].n4 5.02496
R7392 uo_out[6].n4 uo_out[6].n2 0.438
R7393 uo_out[6] uo_out[6].n5 0.063
R7394 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t7 628.097
R7395 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t5 622.766
R7396 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t3 523.774
R7397 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t4 304.647
R7398 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t6 304.647
R7399 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t2 202.44
R7400 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 169.062
R7401 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 166.237
R7402 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t0 84.7557
R7403 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t1 84.1197
R7404 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 12.6535
R7405 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 5.48979
R7406 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 4.5005
R7407 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 1.09595
R7408 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t13 539.841
R7409 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t8 539.841
R7410 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t9 539.841
R7411 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t12 539.841
R7412 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t11 215.293
R7413 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t14 215.293
R7414 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t15 215.293
R7415 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t10 215.293
R7416 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 166.144
R7417 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 165.8
R7418 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t5 85.2499
R7419 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t0 85.2499
R7420 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t3 83.7172
R7421 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t7 83.7172
R7422 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 75.7282
R7423 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 66.3172
R7424 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 36.1505
R7425 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 36.1505
R7426 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 34.5438
R7427 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 34.5438
R7428 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t1 17.4005
R7429 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t2 17.4005
R7430 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t6 9.52217
R7431 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t4 9.52217
R7432 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 6.39571
R7433 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 5.30824
R7434 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 4.94887
R7435 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 1.06691
R7436 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 0.160656
R7437 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t10 539.841
R7438 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t13 539.841
R7439 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t14 539.841
R7440 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t8 539.841
R7441 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t9 215.293
R7442 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t11 215.293
R7443 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t12 215.293
R7444 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t15 215.293
R7445 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 166.149
R7446 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 165.8
R7447 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t2 85.1574
R7448 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t0 85.1574
R7449 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t1 83.8097
R7450 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t7 83.8097
R7451 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 74.288
R7452 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 67.7574
R7453 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 36.1505
R7454 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 36.1505
R7455 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 34.5438
R7456 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 34.5438
R7457 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t3 17.4005
R7458 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t4 17.4005
R7459 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 11.8364
R7460 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t5 9.52217
R7461 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t6 9.52217
R7462 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 5.83219
R7463 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 5.74235
R7464 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 5.49235
R7465 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 1.32081
R7466 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 0.285656
R7467 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t12 539.841
R7468 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t14 539.841
R7469 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t8 539.841
R7470 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t11 539.841
R7471 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t10 215.293
R7472 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t13 215.293
R7473 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t15 215.293
R7474 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t9 215.293
R7475 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 166.144
R7476 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 165.8
R7477 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t6 85.2499
R7478 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t2 85.2499
R7479 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t7 83.7172
R7480 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t3 83.7172
R7481 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 75.7282
R7482 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 66.3172
R7483 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 36.1505
R7484 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 36.1505
R7485 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 34.5438
R7486 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 34.5438
R7487 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t1 17.4005
R7488 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t5 17.4005
R7489 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t4 9.52217
R7490 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t0 9.52217
R7491 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 6.39571
R7492 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 5.30824
R7493 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 4.94887
R7494 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 1.41456
R7495 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t9 539.841
R7496 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t12 539.841
R7497 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t11 539.841
R7498 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t14 539.841
R7499 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t15 215.293
R7500 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t10 215.293
R7501 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t8 215.293
R7502 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t13 215.293
R7503 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 166.149
R7504 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 165.8
R7505 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t0 85.1574
R7506 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t4 85.1574
R7507 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t7 83.8097
R7508 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t1 83.8097
R7509 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 74.288
R7510 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 67.7574
R7511 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 36.1505
R7512 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 36.1505
R7513 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 34.5438
R7514 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 34.5438
R7515 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t5 17.4005
R7516 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t2 17.4005
R7517 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 11.8364
R7518 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t3 9.52217
R7519 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t6 9.52217
R7520 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 5.83219
R7521 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 5.74235
R7522 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 5.49235
R7523 tdc_0.diff_gen_0.delay_unit_2_4.out_1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 1.32081
R7524 tdc_0.diff_gen_0.delay_unit_2_4.out_1 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 0.53175
R7525 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 552.84
R7526 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 552.84
R7527 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 552.84
R7528 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 552.84
R7529 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 539.841
R7530 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 539.841
R7531 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 539.841
R7532 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 539.841
R7533 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 215.293
R7534 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 215.293
R7535 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 215.293
R7536 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 215.293
R7537 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 166.468
R7538 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 166.149
R7539 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 165.8
R7540 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 165.8
R7541 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 85.1574
R7542 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 83.8097
R7543 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 83.8097
R7544 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 83.7172
R7545 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 74.288
R7546 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 67.7574
R7547 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 36.1505
R7548 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 36.1505
R7549 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 34.5438
R7550 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 34.5438
R7551 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 17.4005
R7552 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 17.4005
R7553 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 16.09
R7554 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 11.8364
R7555 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 9.52217
R7556 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 9.52217
R7557 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 5.96628
R7558 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 5.83219
R7559 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 5.74235
R7560 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 5.49235
R7561 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 1.44072
R7562 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 1.32081
R7563 a_10958_34774.n2 a_10958_34774.t3 31.9657
R7564 a_10958_34774.n2 a_10958_34774.n1 25.8125
R7565 a_10958_34774.n4 a_10958_34774.n3 25.8125
R7566 a_10958_34774.n6 a_10958_34774.n5 25.8125
R7567 a_10958_34774.n9 a_10958_34774.n0 25.7038
R7568 a_10958_34774.n10 a_10958_34774.n9 25.3505
R7569 a_10958_34774.n8 a_10958_34774.n7 24.288
R7570 a_10958_34774.n7 a_10958_34774.t7 5.8005
R7571 a_10958_34774.n7 a_10958_34774.t11 5.8005
R7572 a_10958_34774.n1 a_10958_34774.t12 5.8005
R7573 a_10958_34774.n1 a_10958_34774.t0 5.8005
R7574 a_10958_34774.n3 a_10958_34774.t2 5.8005
R7575 a_10958_34774.n3 a_10958_34774.t4 5.8005
R7576 a_10958_34774.n5 a_10958_34774.t10 5.8005
R7577 a_10958_34774.n5 a_10958_34774.t1 5.8005
R7578 a_10958_34774.n0 a_10958_34774.t6 5.8005
R7579 a_10958_34774.n0 a_10958_34774.t8 5.8005
R7580 a_10958_34774.t9 a_10958_34774.n10 5.8005
R7581 a_10958_34774.n10 a_10958_34774.t5 5.8005
R7582 a_10958_34774.n8 a_10958_34774.n6 1.87822
R7583 a_10958_34774.n9 a_10958_34774.n8 1.41626
R7584 a_10958_34774.n4 a_10958_34774.n2 0.353761
R7585 a_10958_34774.n6 a_10958_34774.n4 0.353761
R7586 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t14 539.841
R7587 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t8 539.841
R7588 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t10 539.841
R7589 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t13 539.841
R7590 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t12 215.293
R7591 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t15 215.293
R7592 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t9 215.293
R7593 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t11 215.293
R7594 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 166.144
R7595 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 165.8
R7596 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t5 85.2499
R7597 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t7 85.2499
R7598 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t0 83.7172
R7599 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t6 83.7172
R7600 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 75.7282
R7601 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 66.3172
R7602 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 36.1505
R7603 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 36.1505
R7604 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 34.5438
R7605 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 34.5438
R7606 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t1 17.4005
R7607 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t3 17.4005
R7608 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t4 9.52217
R7609 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t2 9.52217
R7610 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 6.39571
R7611 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 5.30824
R7612 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 4.94887
R7613 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 1.41456
R7614 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 784.053
R7615 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 784.053
R7616 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 784.053
R7617 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 784.053
R7618 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 539.841
R7619 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 539.841
R7620 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 539.841
R7621 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 539.841
R7622 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 215.293
R7623 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 215.293
R7624 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 215.293
R7625 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 215.293
R7626 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 168.659
R7627 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 167.992
R7628 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 166.144
R7629 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 165.8
R7630 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 85.2499
R7631 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 85.2499
R7632 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 83.7172
R7633 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 83.7172
R7634 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 75.7282
R7635 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 66.3172
R7636 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 36.1505
R7637 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 36.1505
R7638 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 34.5438
R7639 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 34.5438
R7640 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 17.4005
R7641 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 17.4005
R7642 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 17.2391
R7643 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 9.52217
R7644 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 9.52217
R7645 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 6.39571
R7646 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 5.30824
R7647 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 4.94887
R7648 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 1.06691
R7649 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 890.727
R7650 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 742.783
R7651 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 641.061
R7652 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 623.388
R7653 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 547.874
R7654 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 431.807
R7655 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 427.875
R7656 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 340.632
R7657 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 208.631
R7658 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 168.007
R7659 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R7660 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 31.2103
R7661 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 31.0962
R7662 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R7663 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R7664 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 8.91506
R7665 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R7666 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R7667 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R7668 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R7669 uo_out[5].n0 uo_out[5].t4 734.539
R7670 uo_out[5].n0 uo_out[5].t5 233.26
R7671 uo_out[5].n2 uo_out[5].n0 162.335
R7672 uo_out[5].n2 uo_out[5].n1 75.5733
R7673 uo_out[5].n4 uo_out[5].n3 66.3172
R7674 uo_out[5].n5 uo_out[5] 19.2682
R7675 uo_out[5].n3 uo_out[5].t1 17.4005
R7676 uo_out[5].n3 uo_out[5].t2 17.4005
R7677 uo_out[5].n1 uo_out[5].t3 9.52217
R7678 uo_out[5].n1 uo_out[5].t0 9.52217
R7679 uo_out[5].n5 uo_out[5].n4 5.02496
R7680 uo_out[5].n4 uo_out[5].n2 0.438
R7681 uo_out[5] uo_out[5].n5 0.063
R7682 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 552.84
R7683 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 552.84
R7684 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 552.84
R7685 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 552.84
R7686 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 539.841
R7687 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 539.841
R7688 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 539.841
R7689 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 539.841
R7690 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 215.293
R7691 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 215.293
R7692 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 215.293
R7693 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 215.293
R7694 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 166.468
R7695 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 166.149
R7696 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 165.8
R7697 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 165.8
R7698 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 85.1574
R7699 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 83.8097
R7700 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 83.8097
R7701 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 83.7172
R7702 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 74.288
R7703 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 67.7574
R7704 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 36.1505
R7705 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 36.1505
R7706 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 34.5438
R7707 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 34.5438
R7708 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 17.4005
R7709 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 17.4005
R7710 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 16.09
R7711 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 11.8364
R7712 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 9.52217
R7713 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 9.52217
R7714 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 5.96628
R7715 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 5.83219
R7716 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 5.74235
R7717 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 5.49235
R7718 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 1.44072
R7719 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 1.32081
R7720 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 0.285656
R7721 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t7 628.097
R7722 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t5 622.766
R7723 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t3 523.774
R7724 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t4 304.647
R7725 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t6 304.647
R7726 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t2 202.44
R7727 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 169.062
R7728 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 166.237
R7729 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t0 84.7557
R7730 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t1 84.1197
R7731 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 12.6535
R7732 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 5.48979
R7733 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 4.5005
R7734 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 1.09595
R7735 ui_in[5].n0 ui_in[5].t7 628.097
R7736 ui_in[5].n1 ui_in[5].t3 622.766
R7737 ui_in[5].n5 ui_in[5].t0 543.053
R7738 ui_in[5].n0 ui_in[5].t5 523.774
R7739 ui_in[5].n2 ui_in[5].t6 304.647
R7740 ui_in[5].n2 ui_in[5].t2 304.647
R7741 ui_in[5].n5 ui_in[5].t1 221.72
R7742 ui_in[5].n6 ui_in[5].n5 220.327
R7743 ui_in[5].n2 ui_in[5].t4 202.44
R7744 ui_in[5] ui_in[5].n2 169.071
R7745 ui_in[5] ui_in[5].n1 166.244
R7746 ui_in[5].n4 ui_in[5] 30.5822
R7747 ui_in[5].n4 ui_in[5].n3 3.0755
R7748 ui_in[5].n3 ui_in[5] 1.24128
R7749 ui_in[5].n1 ui_in[5].n0 1.09595
R7750 ui_in[5].n3 ui_in[5] 0.402286
R7751 ui_in[5].n6 ui_in[5] 0.063
R7752 ui_in[5] ui_in[5].n6 0.0505
R7753 ui_in[5] ui_in[5].n4 0.0147857
R7754 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t9 539.841
R7755 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t11 539.841
R7756 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t13 539.841
R7757 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t8 539.841
R7758 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t15 215.293
R7759 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t10 215.293
R7760 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t12 215.293
R7761 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t14 215.293
R7762 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 166.144
R7763 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 165.8
R7764 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t5 85.2499
R7765 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t1 85.2499
R7766 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t3 83.7172
R7767 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t0 83.7172
R7768 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 75.7282
R7769 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 66.3172
R7770 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 36.1505
R7771 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 36.1505
R7772 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 34.5438
R7773 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 34.5438
R7774 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t4 17.4005
R7775 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t2 17.4005
R7776 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t6 9.52217
R7777 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t7 9.52217
R7778 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 6.39571
R7779 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 5.30824
R7780 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 4.94887
R7781 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 1.06691
R7782 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 0.160656
R7783 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t14 539.841
R7784 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t11 539.841
R7785 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t9 539.841
R7786 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t12 539.841
R7787 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t13 215.293
R7788 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t8 215.293
R7789 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t15 215.293
R7790 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t10 215.293
R7791 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 166.149
R7792 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 165.8
R7793 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t2 85.1574
R7794 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t6 85.1574
R7795 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t3 83.8097
R7796 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t7 83.8097
R7797 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 74.288
R7798 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 67.7574
R7799 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 36.1505
R7800 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 36.1505
R7801 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 34.5438
R7802 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 34.5438
R7803 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t0 17.4005
R7804 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t1 17.4005
R7805 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 11.8364
R7806 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t4 9.52217
R7807 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t5 9.52217
R7808 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 5.83219
R7809 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 5.74235
R7810 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 5.49235
R7811 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 1.32081
R7812 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 0.285656
R7813 a_10958_27928.n2 a_10958_27928.t12 31.9657
R7814 a_10958_27928.n2 a_10958_27928.n1 25.8125
R7815 a_10958_27928.n4 a_10958_27928.n3 25.8125
R7816 a_10958_27928.n6 a_10958_27928.n5 25.8125
R7817 a_10958_27928.n9 a_10958_27928.n0 25.7038
R7818 a_10958_27928.n10 a_10958_27928.n9 25.3505
R7819 a_10958_27928.n8 a_10958_27928.n7 24.288
R7820 a_10958_27928.n7 a_10958_27928.t6 5.8005
R7821 a_10958_27928.n7 a_10958_27928.t1 5.8005
R7822 a_10958_27928.n1 a_10958_27928.t2 5.8005
R7823 a_10958_27928.n1 a_10958_27928.t9 5.8005
R7824 a_10958_27928.n3 a_10958_27928.t11 5.8005
R7825 a_10958_27928.n3 a_10958_27928.t0 5.8005
R7826 a_10958_27928.n5 a_10958_27928.t3 5.8005
R7827 a_10958_27928.n5 a_10958_27928.t10 5.8005
R7828 a_10958_27928.n0 a_10958_27928.t4 5.8005
R7829 a_10958_27928.n0 a_10958_27928.t7 5.8005
R7830 a_10958_27928.t8 a_10958_27928.n10 5.8005
R7831 a_10958_27928.n10 a_10958_27928.t5 5.8005
R7832 a_10958_27928.n8 a_10958_27928.n6 1.87822
R7833 a_10958_27928.n9 a_10958_27928.n8 1.41626
R7834 a_10958_27928.n4 a_10958_27928.n2 0.353761
R7835 a_10958_27928.n6 a_10958_27928.n4 0.353761
R7836 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 879.481
R7837 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 742.783
R7838 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 641.061
R7839 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 623.388
R7840 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 547.874
R7841 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 431.807
R7842 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 427.875
R7843 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 333.161
R7844 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 208.668
R7845 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 168.077
R7846 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 75.5951
R7847 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R7848 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R7849 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 11.1806
R7850 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R7851 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R7852 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R7853 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R7854 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t6 628.097
R7855 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t3 622.766
R7856 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t2 523.774
R7857 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t5 304.647
R7858 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t7 304.647
R7859 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t4 202.44
R7860 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 169.062
R7861 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 166.237
R7862 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t1 84.7557
R7863 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t0 84.1197
R7864 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 12.6535
R7865 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 5.48979
R7866 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en 4.5005
R7867 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 1.09595
R7868 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 784.053
R7869 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 784.053
R7870 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 784.053
R7871 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 784.053
R7872 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 539.841
R7873 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 539.841
R7874 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 539.841
R7875 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 539.841
R7876 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 215.293
R7877 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 215.293
R7878 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 215.293
R7879 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 215.293
R7880 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 168.659
R7881 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 167.992
R7882 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 166.144
R7883 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 165.8
R7884 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 85.2499
R7885 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 85.2499
R7886 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 83.7172
R7887 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 83.7172
R7888 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 75.7282
R7889 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 66.3172
R7890 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 36.1505
R7891 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 36.1505
R7892 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 34.5438
R7893 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 34.5438
R7894 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 17.4005
R7895 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 17.4005
R7896 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 17.2391
R7897 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 9.52217
R7898 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 9.52217
R7899 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 6.39571
R7900 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 5.30824
R7901 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 4.94887
R7902 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 1.06691
R7903 a_10108_30826.n2 a_10108_30826.n1 34.9195
R7904 a_10108_30826.n3 a_10108_30826.n2 25.5407
R7905 a_10108_30826.n2 a_10108_30826.n0 25.2907
R7906 a_10108_30826.n1 a_10108_30826.t3 5.8005
R7907 a_10108_30826.n1 a_10108_30826.t4 5.8005
R7908 a_10108_30826.n0 a_10108_30826.t2 5.8005
R7909 a_10108_30826.n0 a_10108_30826.t5 5.8005
R7910 a_10108_30826.n3 a_10108_30826.t0 5.8005
R7911 a_10108_30826.t1 a_10108_30826.n3 5.8005
R7912 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 784.053
R7913 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 784.053
R7914 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 784.053
R7915 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 784.053
R7916 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 539.841
R7917 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 539.841
R7918 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 539.841
R7919 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 539.841
R7920 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 215.293
R7921 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 215.293
R7922 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 215.293
R7923 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 215.293
R7924 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 168.659
R7925 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 167.992
R7926 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 166.144
R7927 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 165.8
R7928 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 85.2499
R7929 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 85.2499
R7930 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 83.7172
R7931 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 83.7172
R7932 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 75.7282
R7933 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 66.3172
R7934 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 36.1505
R7935 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 36.1505
R7936 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 34.5438
R7937 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 34.5438
R7938 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 17.4005
R7939 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 17.4005
R7940 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 17.2391
R7941 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 9.52217
R7942 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 9.52217
R7943 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 6.39571
R7944 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 5.30824
R7945 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 4.94887
R7946 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 1.06691
R7947 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t13 539.841
R7948 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t8 539.841
R7949 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t9 539.841
R7950 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t11 539.841
R7951 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t12 215.293
R7952 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t14 215.293
R7953 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t15 215.293
R7954 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t10 215.293
R7955 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 166.149
R7956 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 165.8
R7957 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t2 85.1574
R7958 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t0 85.1574
R7959 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t5 83.8097
R7960 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t1 83.8097
R7961 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 74.288
R7962 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 67.7574
R7963 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 36.1505
R7964 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 36.1505
R7965 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 34.5438
R7966 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 34.5438
R7967 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t3 17.4005
R7968 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t4 17.4005
R7969 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 11.8364
R7970 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t6 9.52217
R7971 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t7 9.52217
R7972 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 5.83219
R7973 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 5.74235
R7974 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 5.49235
R7975 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 1.32081
R7976 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 0.285656
R7977 uo_out[0].n0 uo_out[0].t5 734.539
R7978 uo_out[0].n0 uo_out[0].t4 233.26
R7979 uo_out[0].n2 uo_out[0].n0 162.335
R7980 uo_out[0].n2 uo_out[0].n1 75.5733
R7981 uo_out[0].n4 uo_out[0].n3 66.3172
R7982 uo_out[0].n5 uo_out[0] 33.5966
R7983 uo_out[0].n3 uo_out[0].t2 17.4005
R7984 uo_out[0].n3 uo_out[0].t0 17.4005
R7985 uo_out[0].n1 uo_out[0].t1 9.52217
R7986 uo_out[0].n1 uo_out[0].t3 9.52217
R7987 uo_out[0].n5 uo_out[0].n4 5.02496
R7988 uo_out[0].n4 uo_out[0].n2 0.438
R7989 uo_out[0] uo_out[0].n5 0.063
R7990 a_10958_25646.n1 a_10958_25646.t5 31.9657
R7991 a_10958_25646.n1 a_10958_25646.n0 25.8125
R7992 a_10958_25646.n3 a_10958_25646.n2 25.8125
R7993 a_10958_25646.n5 a_10958_25646.n4 25.8125
R7994 a_10958_25646.n10 a_10958_25646.n9 25.7038
R7995 a_10958_25646.n9 a_10958_25646.n8 25.3505
R7996 a_10958_25646.n7 a_10958_25646.n6 24.288
R7997 a_10958_25646.n6 a_10958_25646.t12 5.8005
R7998 a_10958_25646.n6 a_10958_25646.t3 5.8005
R7999 a_10958_25646.n0 a_10958_25646.t2 5.8005
R8000 a_10958_25646.n0 a_10958_25646.t6 5.8005
R8001 a_10958_25646.n2 a_10958_25646.t4 5.8005
R8002 a_10958_25646.n2 a_10958_25646.t1 5.8005
R8003 a_10958_25646.n4 a_10958_25646.t0 5.8005
R8004 a_10958_25646.n4 a_10958_25646.t7 5.8005
R8005 a_10958_25646.n8 a_10958_25646.t8 5.8005
R8006 a_10958_25646.n8 a_10958_25646.t9 5.8005
R8007 a_10958_25646.n10 a_10958_25646.t10 5.8005
R8008 a_10958_25646.t11 a_10958_25646.n10 5.8005
R8009 a_10958_25646.n7 a_10958_25646.n5 1.87822
R8010 a_10958_25646.n9 a_10958_25646.n7 1.41626
R8011 a_10958_25646.n3 a_10958_25646.n1 0.353761
R8012 a_10958_25646.n5 a_10958_25646.n3 0.353761
R8013 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 890.727
R8014 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 742.783
R8015 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 641.061
R8016 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 623.388
R8017 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 547.874
R8018 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 431.807
R8019 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 427.875
R8020 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 340.632
R8021 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 208.631
R8022 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 168.007
R8023 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R8024 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 31.2103
R8025 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 31.0962
R8026 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R8027 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R8028 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 8.91506
R8029 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R8030 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R8031 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R8032 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R8033 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 879.481
R8034 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 742.783
R8035 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 641.061
R8036 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 623.388
R8037 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 547.874
R8038 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 431.807
R8039 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 427.875
R8040 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 333.161
R8041 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 208.668
R8042 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 168.077
R8043 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 75.5951
R8044 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R8045 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R8046 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 11.1806
R8047 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 10.4291
R8048 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R8049 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R8050 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 0.740618
R8051 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 0.228761
R8052 uo_out[3].n0 uo_out[3].t4 734.539
R8053 uo_out[3].n0 uo_out[3].t5 233.26
R8054 uo_out[3].n2 uo_out[3].n0 162.335
R8055 uo_out[3].n2 uo_out[3].n1 75.5733
R8056 uo_out[3].n4 uo_out[3].n3 66.3172
R8057 uo_out[3].n5 uo_out[3] 24.9996
R8058 uo_out[3].n3 uo_out[3].t2 17.4005
R8059 uo_out[3].n3 uo_out[3].t1 17.4005
R8060 uo_out[3].n1 uo_out[3].t0 9.52217
R8061 uo_out[3].n1 uo_out[3].t3 9.52217
R8062 uo_out[3].n5 uo_out[3].n4 5.02496
R8063 uo_out[3].n4 uo_out[3].n2 0.438
R8064 uo_out[3] uo_out[3].n5 0.063
R8065 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t7 628.097
R8066 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t5 622.766
R8067 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t3 523.774
R8068 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t6 304.647
R8069 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t2 304.647
R8070 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t4 202.44
R8071 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 169.062
R8072 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 166.237
R8073 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t1 84.7557
R8074 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t0 84.1197
R8075 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 12.6535
R8076 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 5.48979
R8077 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 4.5005
R8078 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 1.09595
R8079 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t10 539.841
R8080 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t13 539.841
R8081 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t14 539.841
R8082 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t9 539.841
R8083 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t8 215.293
R8084 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t11 215.293
R8085 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t12 215.293
R8086 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t15 215.293
R8087 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 166.144
R8088 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 165.8
R8089 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t3 85.2499
R8090 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t1 85.2499
R8091 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t7 83.7172
R8092 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t2 83.7172
R8093 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 75.7282
R8094 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 66.3172
R8095 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 36.1505
R8096 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 36.1505
R8097 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 34.5438
R8098 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 34.5438
R8099 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t0 17.4005
R8100 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t6 17.4005
R8101 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t4 9.52217
R8102 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t5 9.52217
R8103 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 6.39571
R8104 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 5.30824
R8105 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 4.94887
R8106 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 1.41456
R8107 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t8 539.841
R8108 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t11 539.841
R8109 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t12 539.841
R8110 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t14 539.841
R8111 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t15 215.293
R8112 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t9 215.293
R8113 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t10 215.293
R8114 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t13 215.293
R8115 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 166.149
R8116 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 165.8
R8117 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t1 85.1574
R8118 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t6 85.1574
R8119 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t3 83.8097
R8120 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t7 83.8097
R8121 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 74.288
R8122 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 67.7574
R8123 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 36.1505
R8124 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 36.1505
R8125 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 34.5438
R8126 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 34.5438
R8127 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t2 17.4005
R8128 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t0 17.4005
R8129 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 11.8364
R8130 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t4 9.52217
R8131 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t5 9.52217
R8132 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 5.83219
R8133 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 5.74235
R8134 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 5.49235
R8135 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 1.32081
R8136 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 0.285656
R8137 a_10958_32492.n1 a_10958_32492.t5 31.9657
R8138 a_10958_32492.n1 a_10958_32492.n0 25.8125
R8139 a_10958_32492.n3 a_10958_32492.n2 25.8125
R8140 a_10958_32492.n5 a_10958_32492.n4 25.8125
R8141 a_10958_32492.n10 a_10958_32492.n9 25.7038
R8142 a_10958_32492.n9 a_10958_32492.n8 25.3505
R8143 a_10958_32492.n7 a_10958_32492.n6 24.288
R8144 a_10958_32492.n6 a_10958_32492.t10 5.8005
R8145 a_10958_32492.n6 a_10958_32492.t12 5.8005
R8146 a_10958_32492.n0 a_10958_32492.t4 5.8005
R8147 a_10958_32492.n0 a_10958_32492.t6 5.8005
R8148 a_10958_32492.n2 a_10958_32492.t0 5.8005
R8149 a_10958_32492.n2 a_10958_32492.t3 5.8005
R8150 a_10958_32492.n4 a_10958_32492.t2 5.8005
R8151 a_10958_32492.n4 a_10958_32492.t1 5.8005
R8152 a_10958_32492.n8 a_10958_32492.t8 5.8005
R8153 a_10958_32492.n8 a_10958_32492.t9 5.8005
R8154 a_10958_32492.t11 a_10958_32492.n10 5.8005
R8155 a_10958_32492.n10 a_10958_32492.t7 5.8005
R8156 a_10958_32492.n7 a_10958_32492.n5 1.87822
R8157 a_10958_32492.n9 a_10958_32492.n7 1.41626
R8158 a_10958_32492.n3 a_10958_32492.n1 0.353761
R8159 a_10958_32492.n5 a_10958_32492.n3 0.353761
R8160 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 552.84
R8161 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 552.84
R8162 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 552.84
R8163 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 552.84
R8164 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 539.841
R8165 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 539.841
R8166 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 539.841
R8167 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 539.841
R8168 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 215.293
R8169 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 215.293
R8170 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 215.293
R8171 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 215.293
R8172 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 166.468
R8173 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 166.149
R8174 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 165.8
R8175 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 165.8
R8176 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 85.1574
R8177 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 83.8097
R8178 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 83.8097
R8179 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 83.7172
R8180 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 74.288
R8181 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 67.7574
R8182 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 36.1505
R8183 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 36.1505
R8184 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 34.5438
R8185 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 34.5438
R8186 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 17.4005
R8187 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 17.4005
R8188 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 16.09
R8189 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 11.8364
R8190 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 9.52217
R8191 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 9.52217
R8192 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 5.96628
R8193 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 5.83219
R8194 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 5.74235
R8195 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 5.49235
R8196 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 1.44072
R8197 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 1.32081
R8198 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t13 539.841
R8199 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t9 539.841
R8200 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t8 539.841
R8201 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t11 539.841
R8202 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t12 215.293
R8203 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t15 215.293
R8204 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t14 215.293
R8205 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t10 215.293
R8206 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 166.149
R8207 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 165.8
R8208 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t0 85.1574
R8209 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t6 85.1574
R8210 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t7 83.8097
R8211 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t5 83.8097
R8212 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 74.288
R8213 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 67.7574
R8214 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 36.1505
R8215 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 36.1505
R8216 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 34.5438
R8217 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 34.5438
R8218 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t1 17.4005
R8219 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t2 17.4005
R8220 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 11.8364
R8221 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t3 9.52217
R8222 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t4 9.52217
R8223 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 5.83219
R8224 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 5.74235
R8225 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 5.49235
R8226 tdc_0.diff_gen_0.delay_unit_2_1.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 1.32081
R8227 tdc_0.diff_gen_0.delay_unit_2_1.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 0.285656
R8228 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 784.053
R8229 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 784.053
R8230 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 784.053
R8231 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 784.053
R8232 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 539.841
R8233 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 539.841
R8234 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 539.841
R8235 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 539.841
R8236 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 215.293
R8237 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 215.293
R8238 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 215.293
R8239 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 215.293
R8240 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 168.659
R8241 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 167.992
R8242 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 166.144
R8243 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 165.8
R8244 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 85.2499
R8245 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 85.2499
R8246 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 83.7172
R8247 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 83.7172
R8248 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 75.7282
R8249 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 66.3172
R8250 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 36.1505
R8251 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 36.1505
R8252 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 34.5438
R8253 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 34.5438
R8254 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 17.4005
R8255 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 17.4005
R8256 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 17.2391
R8257 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 9.52217
R8258 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 9.52217
R8259 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 6.39571
R8260 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 5.30824
R8261 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 4.94887
R8262 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 1.06691
R8263 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 879.481
R8264 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 742.783
R8265 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 641.061
R8266 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 623.388
R8267 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 547.874
R8268 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 431.807
R8269 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 427.875
R8270 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 333.161
R8271 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 208.668
R8272 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 168.077
R8273 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 75.5951
R8274 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 31.2972
R8275 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 31.2972
R8276 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 11.1806
R8277 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 10.4291
R8278 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R8279 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R8280 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 0.968879
R8281 variable_delay_short_0.variable_delay_unit_5.in.n0 variable_delay_short_0.variable_delay_unit_5.in.t5 607.409
R8282 variable_delay_short_0.variable_delay_unit_5.in.n2 variable_delay_short_0.variable_delay_unit_5.in.t2 543.053
R8283 variable_delay_short_0.variable_delay_unit_5.in.n0 variable_delay_short_0.variable_delay_unit_5.in.t4 321.423
R8284 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_5.in.n2 221.778
R8285 variable_delay_short_0.variable_delay_unit_5.in.n2 variable_delay_short_0.variable_delay_unit_5.in.t3 221.72
R8286 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_5.in.n0 161.72
R8287 variable_delay_short_0.variable_delay_unit_5.in.n1 variable_delay_short_0.variable_delay_unit_5.in.t0 84.7227
R8288 variable_delay_short_0.variable_delay_unit_5.in.n1 variable_delay_short_0.variable_delay_unit_5.in.t1 84.0867
R8289 variable_delay_short_0.variable_delay_unit_5.in.n3 variable_delay_short_0.variable_delay_unit_5.in 20.0791
R8290 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_5.in.n3 0.851271
R8291 variable_delay_short_0.variable_delay_unit_5.in.n3 variable_delay_short_0.variable_delay_unit_5.in.n1 0.465495
R8292 variable_delay_short_0.variable_delay_unit_5.forward.n0 variable_delay_short_0.variable_delay_unit_5.forward.t3 607.409
R8293 variable_delay_short_0.variable_delay_unit_5.forward.n0 variable_delay_short_0.variable_delay_unit_5.forward.t2 321.423
R8294 variable_delay_short_0.variable_delay_unit_5.forward variable_delay_short_0.variable_delay_unit_5.forward.n0 161.72
R8295 variable_delay_short_0.variable_delay_unit_5.forward.n1 variable_delay_short_0.variable_delay_unit_5.forward.t1 84.7227
R8296 variable_delay_short_0.variable_delay_unit_5.forward.n1 variable_delay_short_0.variable_delay_unit_5.forward.t0 84.0867
R8297 variable_delay_short_0.variable_delay_unit_5.forward.n2 variable_delay_short_0.variable_delay_unit_5.forward 19.7898
R8298 variable_delay_short_0.variable_delay_unit_5.forward variable_delay_short_0.variable_delay_unit_5.forward.n2 0.851271
R8299 variable_delay_short_0.variable_delay_unit_5.forward.n2 variable_delay_short_0.variable_delay_unit_5.forward.n1 0.465495
R8300 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 552.84
R8301 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 552.84
R8302 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 552.84
R8303 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 552.84
R8304 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 539.841
R8305 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 539.841
R8306 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 539.841
R8307 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 539.841
R8308 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 215.293
R8309 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 215.293
R8310 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 215.293
R8311 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 215.293
R8312 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 166.468
R8313 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 166.149
R8314 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 165.8
R8315 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 165.8
R8316 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 85.1574
R8317 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 83.8097
R8318 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 83.8097
R8319 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 83.7172
R8320 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 74.288
R8321 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 67.7574
R8322 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 36.1505
R8323 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 36.1505
R8324 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 34.5438
R8325 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 34.5438
R8326 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 17.4005
R8327 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 17.4005
R8328 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 16.09
R8329 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 11.8364
R8330 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 9.52217
R8331 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 9.52217
R8332 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 5.96628
R8333 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 5.83219
R8334 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 5.74235
R8335 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 5.49235
R8336 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 1.44072
R8337 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 1.32081
R8338 a_10958_30210.n2 a_10958_30210.t12 31.9657
R8339 a_10958_30210.n2 a_10958_30210.n1 25.8125
R8340 a_10958_30210.n4 a_10958_30210.n3 25.8125
R8341 a_10958_30210.n6 a_10958_30210.n5 25.8125
R8342 a_10958_30210.n9 a_10958_30210.n0 25.7038
R8343 a_10958_30210.n10 a_10958_30210.n9 25.3505
R8344 a_10958_30210.n8 a_10958_30210.n7 24.288
R8345 a_10958_30210.n7 a_10958_30210.t1 5.8005
R8346 a_10958_30210.n7 a_10958_30210.t6 5.8005
R8347 a_10958_30210.n1 a_10958_30210.t5 5.8005
R8348 a_10958_30210.n1 a_10958_30210.t9 5.8005
R8349 a_10958_30210.n3 a_10958_30210.t11 5.8005
R8350 a_10958_30210.n3 a_10958_30210.t7 5.8005
R8351 a_10958_30210.n5 a_10958_30210.t8 5.8005
R8352 a_10958_30210.n5 a_10958_30210.t10 5.8005
R8353 a_10958_30210.n0 a_10958_30210.t0 5.8005
R8354 a_10958_30210.n0 a_10958_30210.t2 5.8005
R8355 a_10958_30210.n10 a_10958_30210.t3 5.8005
R8356 a_10958_30210.t4 a_10958_30210.n10 5.8005
R8357 a_10958_30210.n8 a_10958_30210.n6 1.87822
R8358 a_10958_30210.n9 a_10958_30210.n8 1.41626
R8359 a_10958_30210.n4 a_10958_30210.n2 0.353761
R8360 a_10958_30210.n6 a_10958_30210.n4 0.353761
R8361 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 784.053
R8362 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 784.053
R8363 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 784.053
R8364 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 784.053
R8365 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 539.841
R8366 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 539.841
R8367 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 539.841
R8368 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 539.841
R8369 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 215.293
R8370 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 215.293
R8371 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 215.293
R8372 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 215.293
R8373 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 168.659
R8374 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 167.992
R8375 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 166.144
R8376 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 165.8
R8377 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 85.2499
R8378 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 85.2499
R8379 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 83.7172
R8380 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 83.7172
R8381 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 75.7282
R8382 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 66.3172
R8383 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 36.1505
R8384 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 36.1505
R8385 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 34.5438
R8386 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 34.5438
R8387 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 17.4005
R8388 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 17.4005
R8389 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 17.2391
R8390 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 9.52217
R8391 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 9.52217
R8392 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 6.39571
R8393 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 5.30824
R8394 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 4.94887
R8395 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 1.06691
R8396 a_10108_23980.n3 a_10108_23980.n2 34.9195
R8397 a_10108_23980.n2 a_10108_23980.n1 25.5407
R8398 a_10108_23980.n2 a_10108_23980.n0 25.2907
R8399 a_10108_23980.n1 a_10108_23980.t4 5.8005
R8400 a_10108_23980.n1 a_10108_23980.t5 5.8005
R8401 a_10108_23980.n0 a_10108_23980.t0 5.8005
R8402 a_10108_23980.n0 a_10108_23980.t2 5.8005
R8403 a_10108_23980.n3 a_10108_23980.t1 5.8005
R8404 a_10108_23980.t3 a_10108_23980.n3 5.8005
R8405 variable_delay_short_0.variable_delay_unit_3.in.n0 variable_delay_short_0.variable_delay_unit_3.in.t5 607.409
R8406 variable_delay_short_0.variable_delay_unit_3.in.n2 variable_delay_short_0.variable_delay_unit_3.in.t2 543.053
R8407 variable_delay_short_0.variable_delay_unit_3.in.n0 variable_delay_short_0.variable_delay_unit_3.in.t4 321.423
R8408 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_3.in.n2 221.778
R8409 variable_delay_short_0.variable_delay_unit_3.in.n2 variable_delay_short_0.variable_delay_unit_3.in.t3 221.72
R8410 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_3.in.n0 161.72
R8411 variable_delay_short_0.variable_delay_unit_3.in.n1 variable_delay_short_0.variable_delay_unit_3.in.t1 84.7227
R8412 variable_delay_short_0.variable_delay_unit_3.in.n1 variable_delay_short_0.variable_delay_unit_3.in.t0 84.0867
R8413 variable_delay_short_0.variable_delay_unit_3.in.n3 variable_delay_short_0.variable_delay_unit_3.in 20.0791
R8414 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_3.in.n3 0.851271
R8415 variable_delay_short_0.variable_delay_unit_3.in.n3 variable_delay_short_0.variable_delay_unit_3.in.n1 0.465495
R8416 variable_delay_short_0.variable_delay_unit_4.in.n0 variable_delay_short_0.variable_delay_unit_4.in.t5 607.409
R8417 variable_delay_short_0.variable_delay_unit_4.in.n2 variable_delay_short_0.variable_delay_unit_4.in.t2 543.053
R8418 variable_delay_short_0.variable_delay_unit_4.in.n0 variable_delay_short_0.variable_delay_unit_4.in.t4 321.423
R8419 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_4.in.n2 221.778
R8420 variable_delay_short_0.variable_delay_unit_4.in.n2 variable_delay_short_0.variable_delay_unit_4.in.t3 221.72
R8421 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_4.in.n0 161.72
R8422 variable_delay_short_0.variable_delay_unit_4.in.n1 variable_delay_short_0.variable_delay_unit_4.in.t1 84.7227
R8423 variable_delay_short_0.variable_delay_unit_4.in.n1 variable_delay_short_0.variable_delay_unit_4.in.t0 84.0867
R8424 variable_delay_short_0.variable_delay_unit_4.in.n3 variable_delay_short_0.variable_delay_unit_4.in 20.0791
R8425 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_4.in.n3 0.851271
R8426 variable_delay_short_0.variable_delay_unit_4.in.n3 variable_delay_short_0.variable_delay_unit_4.in.n1 0.465495
R8427 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 552.84
R8428 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 552.84
R8429 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 552.84
R8430 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 552.84
R8431 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 539.841
R8432 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 539.841
R8433 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 539.841
R8434 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 539.841
R8435 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 215.293
R8436 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 215.293
R8437 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 215.293
R8438 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 215.293
R8439 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 166.468
R8440 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 166.149
R8441 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 165.8
R8442 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 165.8
R8443 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 85.1574
R8444 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 83.8097
R8445 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 83.8097
R8446 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 83.7172
R8447 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 74.288
R8448 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 67.7574
R8449 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 36.1505
R8450 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 36.1505
R8451 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 34.5438
R8452 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 34.5438
R8453 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 17.4005
R8454 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 17.4005
R8455 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 16.09
R8456 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 11.8364
R8457 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 9.52217
R8458 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 9.52217
R8459 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 5.96628
R8460 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 5.83219
R8461 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 5.74235
R8462 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 5.49235
R8463 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 1.44072
R8464 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 1.32081
R8465 uo_out[4].n0 uo_out[4].t5 734.539
R8466 uo_out[4].n0 uo_out[4].t4 233.26
R8467 uo_out[4].n2 uo_out[4].n0 162.335
R8468 uo_out[4].n2 uo_out[4].n1 75.5733
R8469 uo_out[4].n4 uo_out[4].n3 66.3172
R8470 uo_out[4].n5 uo_out[4] 22.1339
R8471 uo_out[4].n3 uo_out[4].t3 17.4005
R8472 uo_out[4].n3 uo_out[4].t2 17.4005
R8473 uo_out[4].n1 uo_out[4].t1 9.52217
R8474 uo_out[4].n1 uo_out[4].t0 9.52217
R8475 uo_out[4].n5 uo_out[4].n4 5.02496
R8476 uo_out[4].n4 uo_out[4].n2 0.438
R8477 uo_out[4] uo_out[4].n5 0.063
R8478 ui_in[4].n1 ui_in[4].t2 628.097
R8479 ui_in[4].n2 ui_in[4].t6 622.766
R8480 ui_in[4].n0 ui_in[4].t3 543.053
R8481 ui_in[4].n1 ui_in[4].t0 523.774
R8482 ui_in[4].n3 ui_in[4].t1 304.647
R8483 ui_in[4].n3 ui_in[4].t4 304.647
R8484 ui_in[4].n0 ui_in[4].t5 221.72
R8485 ui_in[4].n6 ui_in[4].n0 220.327
R8486 ui_in[4].n3 ui_in[4].t7 202.44
R8487 ui_in[4] ui_in[4].n3 169.071
R8488 ui_in[4] ui_in[4].n2 166.244
R8489 ui_in[4].n5 ui_in[4] 27.1791
R8490 ui_in[4].n5 ui_in[4].n4 2.98979
R8491 ui_in[4].n4 ui_in[4] 1.24128
R8492 ui_in[4].n2 ui_in[4].n1 1.09595
R8493 ui_in[4].n4 ui_in[4] 0.402286
R8494 ui_in[4].n6 ui_in[4].n5 0.1505
R8495 ui_in[4].n6 ui_in[4] 0.063
R8496 ui_in[4] ui_in[4].n6 0.0219286
R8497 uo_out[7].n0 uo_out[7].t5 734.539
R8498 uo_out[7].n0 uo_out[7].t4 233.26
R8499 uo_out[7].n2 uo_out[7].n0 162.335
R8500 uo_out[7].n2 uo_out[7].n1 75.5733
R8501 uo_out[7].n4 uo_out[7].n3 66.3172
R8502 uo_out[7].n3 uo_out[7].t1 17.4005
R8503 uo_out[7].n3 uo_out[7].t3 17.4005
R8504 uo_out[7].n5 uo_out[7] 13.5368
R8505 uo_out[7].n1 uo_out[7].t2 9.52217
R8506 uo_out[7].n1 uo_out[7].t0 9.52217
R8507 uo_out[7].n5 uo_out[7].n4 5.02496
R8508 uo_out[7].n4 uo_out[7].n2 0.438
R8509 uo_out[7] uo_out[7].n5 0.063
R8510 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 552.84
R8511 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 552.84
R8512 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 552.84
R8513 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 552.84
R8514 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 539.841
R8515 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 539.841
R8516 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 539.841
R8517 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 539.841
R8518 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 215.293
R8519 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 215.293
R8520 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 215.293
R8521 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 215.293
R8522 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 166.468
R8523 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 166.149
R8524 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 165.8
R8525 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 165.8
R8526 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 85.1574
R8527 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 83.8097
R8528 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 83.8097
R8529 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 83.7172
R8530 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 74.288
R8531 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 67.7574
R8532 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 36.1505
R8533 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 36.1505
R8534 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 34.5438
R8535 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 34.5438
R8536 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 17.4005
R8537 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 17.4005
R8538 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 16.09
R8539 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 11.8364
R8540 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 9.52217
R8541 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 9.52217
R8542 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 5.96628
R8543 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 5.83219
R8544 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 5.74235
R8545 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 5.49235
R8546 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 1.44072
R8547 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 1.32081
R8548 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 0.285656
R8549 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t13 539.841
R8550 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t8 539.841
R8551 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t9 539.841
R8552 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t12 539.841
R8553 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t11 215.293
R8554 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t14 215.293
R8555 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t15 215.293
R8556 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t10 215.293
R8557 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 166.144
R8558 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 165.8
R8559 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t6 85.2499
R8560 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t1 85.2499
R8561 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t4 83.7172
R8562 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t0 83.7172
R8563 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 75.7282
R8564 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 66.3172
R8565 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 36.1505
R8566 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 36.1505
R8567 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 34.5438
R8568 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 34.5438
R8569 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t2 17.4005
R8570 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t3 17.4005
R8571 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t7 9.52217
R8572 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t5 9.52217
R8573 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 6.39571
R8574 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 5.30824
R8575 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 4.94887
R8576 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 1.06691
R8577 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 0.160656
R8578 tdc_0.vernier_delay_line_0.start_pos.n1 tdc_0.vernier_delay_line_0.start_pos.t8 539.841
R8579 tdc_0.vernier_delay_line_0.start_pos.n0 tdc_0.vernier_delay_line_0.start_pos.t11 539.841
R8580 tdc_0.vernier_delay_line_0.start_pos.n4 tdc_0.vernier_delay_line_0.start_pos.t12 539.841
R8581 tdc_0.vernier_delay_line_0.start_pos.n3 tdc_0.vernier_delay_line_0.start_pos.t14 539.841
R8582 tdc_0.vernier_delay_line_0.start_pos.n1 tdc_0.vernier_delay_line_0.start_pos.t15 215.293
R8583 tdc_0.vernier_delay_line_0.start_pos.n0 tdc_0.vernier_delay_line_0.start_pos.t9 215.293
R8584 tdc_0.vernier_delay_line_0.start_pos.n4 tdc_0.vernier_delay_line_0.start_pos.t10 215.293
R8585 tdc_0.vernier_delay_line_0.start_pos.n3 tdc_0.vernier_delay_line_0.start_pos.t13 215.293
R8586 tdc_0.vernier_delay_line_0.start_pos.n6 tdc_0.vernier_delay_line_0.start_pos.n2 166.149
R8587 tdc_0.vernier_delay_line_0.start_pos.n6 tdc_0.vernier_delay_line_0.start_pos.n5 165.8
R8588 tdc_0.vernier_delay_line_0.start_pos.n12 tdc_0.vernier_delay_line_0.start_pos.t2 85.1574
R8589 tdc_0.vernier_delay_line_0.start_pos.n7 tdc_0.vernier_delay_line_0.start_pos.t0 85.1574
R8590 tdc_0.vernier_delay_line_0.start_pos.n7 tdc_0.vernier_delay_line_0.start_pos.t1 83.8097
R8591 tdc_0.vernier_delay_line_0.start_pos.n12 tdc_0.vernier_delay_line_0.start_pos.t7 83.8097
R8592 tdc_0.vernier_delay_line_0.start_pos.n11 tdc_0.vernier_delay_line_0.start_pos.n10 74.288
R8593 tdc_0.vernier_delay_line_0.start_pos.n11 tdc_0.vernier_delay_line_0.start_pos.n9 67.7574
R8594 tdc_0.vernier_delay_line_0.start_pos.n2 tdc_0.vernier_delay_line_0.start_pos.n1 36.1505
R8595 tdc_0.vernier_delay_line_0.start_pos.n5 tdc_0.vernier_delay_line_0.start_pos.n3 36.1505
R8596 tdc_0.vernier_delay_line_0.start_pos.n2 tdc_0.vernier_delay_line_0.start_pos.n0 34.5438
R8597 tdc_0.vernier_delay_line_0.start_pos.n5 tdc_0.vernier_delay_line_0.start_pos.n4 34.5438
R8598 tdc_0.vernier_delay_line_0.start_pos.n9 tdc_0.vernier_delay_line_0.start_pos.t3 17.4005
R8599 tdc_0.vernier_delay_line_0.start_pos.n9 tdc_0.vernier_delay_line_0.start_pos.t4 17.4005
R8600 tdc_0.vernier_delay_line_0.start_pos.n8 tdc_0.vernier_delay_line_0.start_pos.n6 11.8364
R8601 tdc_0.vernier_delay_line_0.start_pos.n10 tdc_0.vernier_delay_line_0.start_pos.t5 9.52217
R8602 tdc_0.vernier_delay_line_0.start_pos.n10 tdc_0.vernier_delay_line_0.start_pos.t6 9.52217
R8603 tdc_0.vernier_delay_line_0.start_pos.n13 tdc_0.vernier_delay_line_0.start_pos.n11 5.83219
R8604 tdc_0.vernier_delay_line_0.start_pos.n8 tdc_0.vernier_delay_line_0.start_pos.n7 5.74235
R8605 tdc_0.vernier_delay_line_0.start_pos.n13 tdc_0.vernier_delay_line_0.start_pos.n12 5.49235
R8606 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.start_pos.n13 1.32081
R8607 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.start_pos.n8 0.40675
R8608 ui_in[7].n0 ui_in[7].t5 628.097
R8609 ui_in[7].n1 ui_in[7].t7 622.766
R8610 ui_in[7].n5 ui_in[7].t2 543.053
R8611 ui_in[7].n0 ui_in[7].t1 523.774
R8612 ui_in[7].n2 ui_in[7].t4 304.647
R8613 ui_in[7].n2 ui_in[7].t6 304.647
R8614 ui_in[7].n5 ui_in[7].t3 221.72
R8615 ui_in[7].n6 ui_in[7].n5 220.327
R8616 ui_in[7].n2 ui_in[7].t0 202.44
R8617 ui_in[7] ui_in[7].n2 169.071
R8618 ui_in[7] ui_in[7].n1 166.244
R8619 ui_in[7].n4 ui_in[7] 35.9653
R8620 ui_in[7].n4 ui_in[7].n3 3.04693
R8621 ui_in[7].n3 ui_in[7] 1.24128
R8622 ui_in[7].n1 ui_in[7].n0 1.09595
R8623 ui_in[7].n3 ui_in[7] 0.402286
R8624 ui_in[7].n6 ui_in[7] 0.063
R8625 ui_in[7] ui_in[7].n4 0.0505
R8626 ui_in[7] ui_in[7].n6 0.0433571
R8627 ui_in[6].n0 ui_in[6].t1 628.097
R8628 ui_in[6].n1 ui_in[6].t5 622.766
R8629 ui_in[6].n5 ui_in[6].t2 543.053
R8630 ui_in[6].n0 ui_in[6].t0 523.774
R8631 ui_in[6].n2 ui_in[6].t7 304.647
R8632 ui_in[6].n2 ui_in[6].t4 304.647
R8633 ui_in[6].n5 ui_in[6].t3 221.72
R8634 ui_in[6].n6 ui_in[6].n5 220.327
R8635 ui_in[6].n2 ui_in[6].t6 202.44
R8636 ui_in[6] ui_in[6].n2 169.071
R8637 ui_in[6] ui_in[6].n1 166.244
R8638 ui_in[6].n4 ui_in[6] 33.1777
R8639 ui_in[6].n4 ui_in[6].n3 2.26836
R8640 ui_in[6].n3 ui_in[6] 1.24128
R8641 ui_in[6].n1 ui_in[6].n0 1.09595
R8642 ui_in[6] ui_in[6].n4 0.761214
R8643 ui_in[6].n3 ui_in[6] 0.402286
R8644 ui_in[6] ui_in[6].n6 0.111214
R8645 ui_in[6].n6 ui_in[6] 0.063
R8646 ua[0].n1 ua[0].t2 618.668
R8647 ua[0].n0 ua[0].t3 618.668
R8648 ua[0].n1 ua[0].t0 456.997
R8649 ua[0].n0 ua[0].t1 456.997
R8650 ua[0] ua[0].n1 161.375
R8651 ua[0] ua[0].n0 161.375
R8652 ua[0] ua[0].n2 11.6385
R8653 ua[0].n2 ua[0] 10.7183
R8654 ua[0].n2 ua[0] 5.67014
R8655 uio_in[0].n0 uio_in[0].t5 628.097
R8656 uio_in[0].n1 uio_in[0].t7 622.766
R8657 uio_in[0].n5 uio_in[0].t3 543.053
R8658 uio_in[0].n0 uio_in[0].t1 523.774
R8659 uio_in[0].n2 uio_in[0].t2 304.647
R8660 uio_in[0].n2 uio_in[0].t6 304.647
R8661 uio_in[0].n5 uio_in[0].t4 221.72
R8662 uio_in[0].n6 uio_in[0].n5 220.327
R8663 uio_in[0].n2 uio_in[0].t0 202.44
R8664 uio_in[0] uio_in[0].n2 169.071
R8665 uio_in[0] uio_in[0].n1 166.244
R8666 uio_in[0].n4 uio_in[0] 38.2949
R8667 uio_in[0].n4 uio_in[0].n3 3.06836
R8668 uio_in[0].n3 uio_in[0] 1.24128
R8669 uio_in[0].n1 uio_in[0].n0 1.09595
R8670 uio_in[0].n3 uio_in[0] 0.402286
R8671 uio_in[0].n6 uio_in[0] 0.063
R8672 uio_in[0] uio_in[0].n4 0.0469286
R8673 uio_in[0] uio_in[0].n6 0.0255
R8674 tdc_0.vernier_delay_line_0.start_neg.n2 tdc_0.vernier_delay_line_0.start_neg.t14 539.841
R8675 tdc_0.vernier_delay_line_0.start_neg.n1 tdc_0.vernier_delay_line_0.start_neg.t8 539.841
R8676 tdc_0.vernier_delay_line_0.start_neg.n5 tdc_0.vernier_delay_line_0.start_neg.t11 539.841
R8677 tdc_0.vernier_delay_line_0.start_neg.n4 tdc_0.vernier_delay_line_0.start_neg.t12 539.841
R8678 tdc_0.vernier_delay_line_0.start_neg.n2 tdc_0.vernier_delay_line_0.start_neg.t13 215.293
R8679 tdc_0.vernier_delay_line_0.start_neg.n1 tdc_0.vernier_delay_line_0.start_neg.t15 215.293
R8680 tdc_0.vernier_delay_line_0.start_neg.n5 tdc_0.vernier_delay_line_0.start_neg.t9 215.293
R8681 tdc_0.vernier_delay_line_0.start_neg.n4 tdc_0.vernier_delay_line_0.start_neg.t10 215.293
R8682 tdc_0.vernier_delay_line_0.start_neg.n7 tdc_0.vernier_delay_line_0.start_neg.n3 166.144
R8683 tdc_0.vernier_delay_line_0.start_neg.n7 tdc_0.vernier_delay_line_0.start_neg.n6 165.8
R8684 tdc_0.vernier_delay_line_0.start_neg.n0 tdc_0.vernier_delay_line_0.start_neg.t7 85.2499
R8685 tdc_0.vernier_delay_line_0.start_neg.n11 tdc_0.vernier_delay_line_0.start_neg.t5 85.2499
R8686 tdc_0.vernier_delay_line_0.start_neg.n11 tdc_0.vernier_delay_line_0.start_neg.t0 83.7172
R8687 tdc_0.vernier_delay_line_0.start_neg.n0 tdc_0.vernier_delay_line_0.start_neg.t6 83.7172
R8688 tdc_0.vernier_delay_line_0.start_neg.n10 tdc_0.vernier_delay_line_0.start_neg.n8 75.7282
R8689 tdc_0.vernier_delay_line_0.start_neg.n10 tdc_0.vernier_delay_line_0.start_neg.n9 66.3172
R8690 tdc_0.vernier_delay_line_0.start_neg.n3 tdc_0.vernier_delay_line_0.start_neg.n1 36.1505
R8691 tdc_0.vernier_delay_line_0.start_neg.n6 tdc_0.vernier_delay_line_0.start_neg.n4 36.1505
R8692 tdc_0.vernier_delay_line_0.start_neg.n3 tdc_0.vernier_delay_line_0.start_neg.n2 34.5438
R8693 tdc_0.vernier_delay_line_0.start_neg.n6 tdc_0.vernier_delay_line_0.start_neg.n5 34.5438
R8694 tdc_0.vernier_delay_line_0.start_neg.n9 tdc_0.vernier_delay_line_0.start_neg.t1 17.4005
R8695 tdc_0.vernier_delay_line_0.start_neg.n9 tdc_0.vernier_delay_line_0.start_neg.t2 17.4005
R8696 tdc_0.vernier_delay_line_0.start_neg.n8 tdc_0.vernier_delay_line_0.start_neg.t3 9.52217
R8697 tdc_0.vernier_delay_line_0.start_neg.n8 tdc_0.vernier_delay_line_0.start_neg.t4 9.52217
R8698 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.start_neg.n0 6.45821
R8699 tdc_0.vernier_delay_line_0.start_neg.n12 tdc_0.vernier_delay_line_0.start_neg.n10 5.30824
R8700 tdc_0.vernier_delay_line_0.start_neg.n12 tdc_0.vernier_delay_line_0.start_neg.n11 4.94887
R8701 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.start_neg.n7 0.754406
R8702 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.start_neg.n12 0.160656
R8703 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 784.053
R8704 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 784.053
R8705 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 784.053
R8706 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 784.053
R8707 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 539.841
R8708 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 539.841
R8709 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 539.841
R8710 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 539.841
R8711 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 215.293
R8712 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 215.293
R8713 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 215.293
R8714 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 215.293
R8715 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 168.659
R8716 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 167.992
R8717 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 166.144
R8718 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 165.8
R8719 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 85.2499
R8720 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 85.2499
R8721 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 83.7172
R8722 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 83.7172
R8723 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 75.7282
R8724 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 66.3172
R8725 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 36.1505
R8726 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 36.1505
R8727 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 34.5438
R8728 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 34.5438
R8729 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 17.4005
R8730 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 17.4005
R8731 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 17.2391
R8732 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 9.52217
R8733 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 9.52217
R8734 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 6.39571
R8735 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 5.30824
R8736 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 4.94887
R8737 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 1.48097
R8738 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 1.06691
R8739 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.539562
R8740 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.391125
R8741 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 0.160656
R8742 a_10108_33108.n3 a_10108_33108.n2 34.9195
R8743 a_10108_33108.n2 a_10108_33108.n1 25.5407
R8744 a_10108_33108.n2 a_10108_33108.n0 25.2907
R8745 a_10108_33108.n1 a_10108_33108.t5 5.8005
R8746 a_10108_33108.n1 a_10108_33108.t4 5.8005
R8747 a_10108_33108.n0 a_10108_33108.t0 5.8005
R8748 a_10108_33108.n0 a_10108_33108.t2 5.8005
R8749 a_10108_33108.n3 a_10108_33108.t1 5.8005
R8750 a_10108_33108.t3 a_10108_33108.n3 5.8005
R8751 variable_delay_dummy_0.variable_delay_unit_1.in.n0 variable_delay_dummy_0.variable_delay_unit_1.in.t4 607.409
R8752 variable_delay_dummy_0.variable_delay_unit_1.in.n2 variable_delay_dummy_0.variable_delay_unit_1.in.t3 543.053
R8753 variable_delay_dummy_0.variable_delay_unit_1.in.n0 variable_delay_dummy_0.variable_delay_unit_1.in.t5 321.423
R8754 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_1.in.n2 221.778
R8755 variable_delay_dummy_0.variable_delay_unit_1.in.n2 variable_delay_dummy_0.variable_delay_unit_1.in.t2 221.72
R8756 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_1.in.n0 161.72
R8757 variable_delay_dummy_0.variable_delay_unit_1.in.n1 variable_delay_dummy_0.variable_delay_unit_1.in.t1 84.7227
R8758 variable_delay_dummy_0.variable_delay_unit_1.in.n1 variable_delay_dummy_0.variable_delay_unit_1.in.t0 84.0867
R8759 variable_delay_dummy_0.variable_delay_unit_1.in.n3 variable_delay_dummy_0.variable_delay_unit_1.in 20.0791
R8760 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_1.in.n3 0.851271
R8761 variable_delay_dummy_0.variable_delay_unit_1.in.n3 variable_delay_dummy_0.variable_delay_unit_1.in.n1 0.465495
R8762 variable_delay_dummy_0.variable_delay_unit_1.forward.n0 variable_delay_dummy_0.variable_delay_unit_1.forward.t2 607.409
R8763 variable_delay_dummy_0.variable_delay_unit_1.forward.n0 variable_delay_dummy_0.variable_delay_unit_1.forward.t3 321.423
R8764 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_1.forward.n0 161.72
R8765 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 variable_delay_dummy_0.variable_delay_unit_1.forward.t1 84.7227
R8766 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 variable_delay_dummy_0.variable_delay_unit_1.forward.t0 84.0867
R8767 variable_delay_dummy_0.variable_delay_unit_1.forward.n2 variable_delay_dummy_0.variable_delay_unit_1.forward 19.7898
R8768 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_1.forward.n2 0.851271
R8769 variable_delay_dummy_0.variable_delay_unit_1.forward.n2 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 0.465495
R8770 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t1 85.1574
R8771 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t3 83.8097
R8772 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 74.288
R8773 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 67.7574
R8774 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t2 17.4005
R8775 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t0 17.4005
R8776 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t4 9.52217
R8777 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t5 9.52217
R8778 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 5.83219
R8779 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 5.49235
R8780 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 1.32081
R8781 ui_in[2].n0 ui_in[2].t0 577.653
R8782 ui_in[2].n0 ui_in[2] 37.1928
R8783 ui_in[2] ui_in[2].n0 0.0747188
R8784 uo_out[1].n0 uo_out[1].t4 734.539
R8785 uo_out[1].n0 uo_out[1].t5 233.26
R8786 uo_out[1].n2 uo_out[1].n0 162.335
R8787 uo_out[1].n2 uo_out[1].n1 75.5733
R8788 uo_out[1].n4 uo_out[1].n3 66.3172
R8789 uo_out[1].n5 uo_out[1] 30.7309
R8790 uo_out[1].n3 uo_out[1].t2 17.4005
R8791 uo_out[1].n3 uo_out[1].t1 17.4005
R8792 uo_out[1].n1 uo_out[1].t0 9.52217
R8793 uo_out[1].n1 uo_out[1].t3 9.52217
R8794 uo_out[1].n5 uo_out[1].n4 5.02496
R8795 uo_out[1].n4 uo_out[1].n2 0.438
R8796 uo_out[1] uo_out[1].n5 0.063
R8797 uo_out[2].n0 uo_out[2].t4 734.539
R8798 uo_out[2].n0 uo_out[2].t5 233.26
R8799 uo_out[2].n2 uo_out[2].n0 162.335
R8800 uo_out[2].n2 uo_out[2].n1 75.5733
R8801 uo_out[2].n4 uo_out[2].n3 66.3172
R8802 uo_out[2].n5 uo_out[2] 27.8652
R8803 uo_out[2].n3 uo_out[2].t0 17.4005
R8804 uo_out[2].n3 uo_out[2].t3 17.4005
R8805 uo_out[2].n1 uo_out[2].t2 9.52217
R8806 uo_out[2].n1 uo_out[2].t1 9.52217
R8807 uo_out[2].n5 uo_out[2].n4 5.02496
R8808 uo_out[2].n4 uo_out[2].n2 0.438
R8809 uo_out[2] uo_out[2].n5 0.063
R8810 uio_in[3].n0 uio_in[3].t0 577.653
R8811 uio_in[3].n0 uio_in[3] 39.6907
R8812 uio_in[3] uio_in[3].n0 0.0747188
R8813 ui_in[0].n0 ui_in[0].t0 577.653
R8814 ui_in[0].n0 ui_in[0] 40.4285
R8815 ui_in[0] ui_in[0].n0 0.0747188
R8816 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 890.727
R8817 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 742.783
R8818 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 641.061
R8819 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 623.388
R8820 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 547.874
R8821 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 431.807
R8822 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 427.875
R8823 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 340.632
R8824 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 208.631
R8825 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 168.007
R8826 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 75.2663
R8827 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 31.2103
R8828 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 31.0962
R8829 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R8830 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R8831 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 8.91506
R8832 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R8833 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R8834 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R8835 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 0.644522
R8836 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 879.481
R8837 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 742.783
R8838 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 641.061
R8839 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 623.388
R8840 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 547.874
R8841 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 431.807
R8842 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 427.875
R8843 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 333.161
R8844 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 208.668
R8845 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 168.077
R8846 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 75.5951
R8847 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 31.2972
R8848 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 31.2972
R8849 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 11.1806
R8850 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 10.4291
R8851 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R8852 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R8853 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 0.740618
R8854 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 0.228761
R8855 a_10108_37672.n3 a_10108_37672.n2 34.9195
R8856 a_10108_37672.n2 a_10108_37672.n1 25.5407
R8857 a_10108_37672.n2 a_10108_37672.n0 25.2907
R8858 a_10108_37672.n1 a_10108_37672.t0 5.8005
R8859 a_10108_37672.n1 a_10108_37672.t1 5.8005
R8860 a_10108_37672.n0 a_10108_37672.t2 5.8005
R8861 a_10108_37672.n0 a_10108_37672.t5 5.8005
R8862 a_10108_37672.n3 a_10108_37672.t3 5.8005
R8863 a_10108_37672.t4 a_10108_37672.n3 5.8005
R8864 variable_delay_short_0.variable_delay_unit_2.in.n0 variable_delay_short_0.variable_delay_unit_2.in.t5 607.409
R8865 variable_delay_short_0.variable_delay_unit_2.in.n2 variable_delay_short_0.variable_delay_unit_2.in.t2 543.053
R8866 variable_delay_short_0.variable_delay_unit_2.in.n0 variable_delay_short_0.variable_delay_unit_2.in.t4 321.423
R8867 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_2.in.n2 221.778
R8868 variable_delay_short_0.variable_delay_unit_2.in.n2 variable_delay_short_0.variable_delay_unit_2.in.t3 221.72
R8869 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_2.in.n0 161.72
R8870 variable_delay_short_0.variable_delay_unit_2.in.n1 variable_delay_short_0.variable_delay_unit_2.in.t0 84.7227
R8871 variable_delay_short_0.variable_delay_unit_2.in.n1 variable_delay_short_0.variable_delay_unit_2.in.t1 84.0867
R8872 variable_delay_short_0.variable_delay_unit_2.in.n3 variable_delay_short_0.variable_delay_unit_2.in 20.0791
R8873 variable_delay_short_0.variable_delay_unit_2.in variable_delay_short_0.variable_delay_unit_2.in.n3 0.851271
R8874 variable_delay_short_0.variable_delay_unit_2.in.n3 variable_delay_short_0.variable_delay_unit_2.in.n1 0.465495
R8875 variable_delay_short_0.variable_delay_unit_1.in.n0 variable_delay_short_0.variable_delay_unit_1.in.t5 607.409
R8876 variable_delay_short_0.variable_delay_unit_1.in.n2 variable_delay_short_0.variable_delay_unit_1.in.t2 543.053
R8877 variable_delay_short_0.variable_delay_unit_1.in.n0 variable_delay_short_0.variable_delay_unit_1.in.t4 321.423
R8878 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_1.in.n2 221.778
R8879 variable_delay_short_0.variable_delay_unit_1.in.n2 variable_delay_short_0.variable_delay_unit_1.in.t3 221.72
R8880 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_1.in.n0 161.72
R8881 variable_delay_short_0.variable_delay_unit_1.in.n1 variable_delay_short_0.variable_delay_unit_1.in.t1 84.7227
R8882 variable_delay_short_0.variable_delay_unit_1.in.n1 variable_delay_short_0.variable_delay_unit_1.in.t0 84.0867
R8883 variable_delay_short_0.variable_delay_unit_1.in.n3 variable_delay_short_0.variable_delay_unit_1.in 20.0791
R8884 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_1.in.n3 0.851271
R8885 variable_delay_short_0.variable_delay_unit_1.in.n3 variable_delay_short_0.variable_delay_unit_1.in.n1 0.465495
R8886 ui_in[3].n0 ui_in[3].t0 727.072
R8887 ui_in[3].n0 ui_in[3] 36.9161
R8888 ui_in[3].n0 ui_in[3] 0.323417
R8889 ui_in[3] ui_in[3].n0 0.0610469
R8890 uio_in[1].n0 uio_in[1].t0 577.653
R8891 uio_in[1].n0 uio_in[1] 42.0234
R8892 uio_in[1] uio_in[1].n0 0.0747188
R8893 uio_in[4].n0 uio_in[4].t0 727.072
R8894 uio_in[4].n0 uio_in[4] 39.7322
R8895 uio_in[4].n0 uio_in[4] 0.323417
R8896 uio_in[4] uio_in[4].n0 0.0610469
R8897 uio_in[5].n0 uio_in[5].t1 564.04
R8898 uio_in[5].n0 uio_in[5].t0 511.623
R8899 uio_in[5].n1 uio_in[5].n0 161.3
R8900 uio_in[5].n1 uio_in[5] 50.8219
R8901 uio_in[5] uio_in[5].n1 0.0295179
R8902 ui_in[1].n0 ui_in[1].t0 727.072
R8903 ui_in[1].n0 ui_in[1] 40.1518
R8904 ui_in[1].n0 ui_in[1] 0.323417
R8905 ui_in[1] ui_in[1].n0 0.0610469
R8906 uio_in[2].n0 uio_in[2].t0 727.072
R8907 uio_in[2].n0 uio_in[2] 42.3292
R8908 uio_in[2].n0 uio_in[2] 0.323417
R8909 uio_in[2] uio_in[2].n0 0.0610469
C0 variable_delay_short_0.variable_delay_unit_1.out ui_in[1] 0.001119f
C1 uio_in[4] variable_delay_dummy_0.in 0.03818f
C2 a_12420_40104# a_12308_40142# 0.030083f
C3 variable_delay_short_0.out tdc_0.diff_gen_0.delay_unit_2_1.in_1 7.3e-20
C4 tdc_0.vernier_delay_line_0.start_neg tdc_0.diff_gen_0.delay_unit_2_6.in_1 0.286409f
C5 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12420_30598# 0.003664f
C6 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12420_37822# 0.003607f
C7 ui_in[6] ui_in[2] 7.13e-19
C8 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12310_32834# 0.014814f
C9 ui_in[4] variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 9.38e-20
C10 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 a_12310_30552# 4.55e-19
C11 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en VDPWR 2.78173f
C12 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 2.36e-21
C13 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_24240_26988# 0.029284f
C14 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.out 0.002141f
C15 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.out 0.235655f
C16 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C17 a_24790_8314# variable_delay_short_0.in 7.3e-20
C18 a_15322_8490# a_16292_8344# 0.019821f
C19 variable_delay_short_0.in VDPWR 1.34358f
C20 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C21 a_12420_26034# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.003664f
C22 variable_delay_dummy_0.in input_stage_0.fine_delay_unit_1.in 0.002924f
C23 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.003768f
C24 uio_out[4] uio_out[3] 0.170937f
C25 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.499806f
C26 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_10108_34862# 0.09966f
C27 a_24240_18144# VDPWR 1.6584f
C28 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 1.99e-19
C29 a_24790_6936# ui_in[1] 0.024305f
C30 a_24240_18144# a_25060_18144# 0.011184f
C31 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.019931f
C32 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.138497f
C33 uio_oe[0] uio_out[7] 0.170937f
C34 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_12308_31014# 7.19e-22
C35 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.99e-19
C36 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en VDPWR 2.7762f
C37 uo_out[3] a_12308_28732# 6.49e-20
C38 a_25060_26988# VDPWR 0.003377f
C39 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12308_33296# 3.26e-19
C40 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_13254_24130# 0.012202f
C41 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 8.54e-19
C42 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 VDPWR 3.23832f
C43 ui_in[7] variable_delay_short_0.variable_delay_unit_2.in 0.574722f
C44 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.out 0.12029f
C45 uio_in[4] a_15322_8490# 0.010812f
C46 uio_in[3] a_16500_11634# 4.35e-20
C47 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_10108_23452# 1.06381f
C48 ui_in[2] variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 6.97e-19
C49 a_12420_39726# VDPWR 0.497771f
C50 uo_out[0] tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.20241f
C51 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.132512f
C52 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 0.085059f
C53 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.441213f
C54 a_16500_12516# variable_delay_dummy_0.in 7.65e-21
C55 a_25060_26988# variable_delay_short_0.variable_delay_unit_5.out 0.172055f
C56 uo_out[0] tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.229249f
C57 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.006183f
C58 ui_in[3] variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.014554f
C59 a_25284_5108# ua[0] 0.009499f
C60 a_23820_8460# a_24790_8314# 0.019821f
C61 a_23820_8460# VDPWR 1.25074f
C62 input_stage_1.fine_delay_unit_0.in ui_in[1] 0.021403f
C63 input_stage_1.fine_delay_unit_1.in variable_delay_short_0.in 0.002949f
C64 a_15322_8490# input_stage_0.fine_delay_unit_1.in 0.254332f
C65 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.003768f
C66 a_12310_35116# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 4.55e-19
C67 a_12310_30552# a_13254_30598# 1.02e-19
C68 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_13254_26412# 0.174293f
C69 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VDPWR 1.93357f
C70 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 a_12310_23706# 4.55e-19
C71 uio_in[4] VDPWR 0.004419f
C72 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.019931f
C73 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.138497f
C74 a_12420_39726# a_12310_39680# 0.030392f
C75 uo_out[1] tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 6.28e-22
C76 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.010157f
C77 a_25060_15196# ui_in[7] 0.001909f
C78 a_16292_8344# a_16292_8080# 0.556904f
C79 variable_delay_short_0.variable_delay_unit_3.in a_24240_18144# 0.020173f
C80 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12310_35116# 0.014814f
C81 ui_in[3] a_25060_12248# 0.002391f
C82 ui_in[5] variable_delay_short_0.variable_delay_unit_4.out 0.043597f
C83 ui_in[5] variable_delay_short_0.variable_delay_unit_5.in 0.00265f
C84 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 7.19e-22
C85 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12308_37860# 2.36e-21
C86 a_12420_39726# uo_out[7] 0.492009f
C87 a_24240_24040# variable_delay_short_0.variable_delay_unit_4.out 0.493816f
C88 a_24240_26106# variable_delay_short_0.variable_delay_unit_5.in 8.82e-20
C89 variable_delay_short_0.variable_delay_unit_5.in a_24240_24040# 0.020173f
C90 input_stage_0.fine_delay_unit_1.in VDPWR 1.33446f
C91 a_13254_30598# VDPWR 6.18e-19
C92 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12310_28270# 0.196592f
C93 variable_delay_short_0.variable_delay_unit_1.in VDPWR 2.13093f
C94 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en VDPWR 3.86957f
C95 a_23820_8460# input_stage_1.fine_delay_unit_1.in 0.254332f
C96 input_stage_1.nand_gate_0.out ui_in[1] 6.37e-19
C97 ui_in[6] a_24240_18144# 0.124274f
C98 uio_in[4] a_16292_8080# 0.00799f
C99 uio_in[5] variable_delay_dummy_0.in 0.060059f
C100 a_12308_35578# uo_out[5] 0.014835f
C101 uio_in[2] a_16292_8344# 4.3e-19
C102 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 9.61e-20
C103 a_15680_15464# variable_delay_dummy_0.variable_delay_unit_1.out 0.493816f
C104 a_13254_40104# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.174293f
C105 uio_in[3] variable_delay_dummy_0.variable_delay_unit_1.in 3.5e-20
C106 a_12310_39680# a_10108_39426# 2.08e-21
C107 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.441213f
C108 a_25060_26106# ui_in[3] 0.002391f
C109 ui_in[3] a_25060_24040# 0.002391f
C110 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.53e-19
C111 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_2 0.667766f
C112 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12420_37444# 0.035356f
C113 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.out 0.12029f
C114 ui_in[6] variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 2.92e-19
C115 ui_in[2] variable_delay_short_0.out 0.003069f
C116 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.in 0.09141f
C117 a_24790_8314# a_24790_8050# 0.556904f
C118 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C119 uo_out[4] VDPWR 0.587468f
C120 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_25060_14314# 2.39e-19
C121 input_stage_0.fine_delay_unit_1.in a_16292_8080# 0.244525f
C122 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.231672f
C123 a_16500_12516# VDPWR 0.003447f
C124 uio_in[4] uio_in[2] 0.01853f
C125 variable_delay_short_0.variable_delay_unit_2.out VDPWR 1.34424f
C126 a_15680_12516# a_16500_12516# 0.011184f
C127 a_25060_18144# variable_delay_short_0.variable_delay_unit_2.out 0.172055f
C128 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 VDPWR 2.23953f
C129 a_12308_24168# a_12420_24130# 0.030083f
C130 variable_delay_short_0.out a_25060_11366# 0.222585f
C131 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 1.99e-19
C132 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 uo_out[4] 1.53e-22
C133 uo_out[0] a_13254_24130# 0.005542f
C134 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 4.28924f
C135 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_12310_23706# 0.164402f
C136 uio_in[5] a_15322_8490# 0.01196f
C137 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.132512f
C138 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 9.61e-20
C139 uio_in[2] input_stage_0.fine_delay_unit_1.in 0.039331f
C140 variable_delay_short_0.variable_delay_unit_1.out ui_in[2] 0.002549f
C141 uio_in[0] VDPWR 1.46811f
C142 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.132512f
C143 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.085059f
C144 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12310_37398# 1.15e-21
C145 a_13254_39726# VDPWR 6.18e-19
C146 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 uo_out[6] 0.20241f
C147 a_16500_14582# VDPWR 0.160518f
C148 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 0.002365f
C149 uio_oe[5] uio_oe[4] 0.170937f
C150 variable_delay_dummy_0.out a_16292_8344# 5.64e-19
C151 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.441213f
C152 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq uo_out[3] 0.229249f
C153 a_25060_20210# VDPWR 6.98e-19
C154 ui_in[3] a_24240_23158# 0.001719f
C155 a_24240_14314# ui_in[7] 0.042718f
C156 input_stage_1.fine_delay_unit_1.in a_24790_8050# 0.244525f
C157 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 1.17e-19
C158 ui_in[7] uio_in[1] 5.13e-19
C159 uo_out[6] uo_out[5] 1.21073f
C160 uo_out[7] uo_out[4] 2.26e-21
C161 tdc_0.vernier_delay_line_0.start_pos VDPWR 4.78299f
C162 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12310_25988# 0.014814f
C163 uio_in[5] VDPWR 0.925517f
C164 uio_in[5] a_15680_12516# 0.002316f
C165 uio_in[4] variable_delay_dummy_0.out 0.007407f
C166 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12308_24168# 7.19e-22
C167 tdc_0.diff_gen_0.delay_unit_2_6.in_2 VDPWR 3.06151f
C168 a_25060_17262# VDPWR 6.98e-19
C169 a_12310_39680# a_13254_39726# 1.02e-19
C170 ui_in[6] variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 2.92e-19
C171 variable_delay_short_0.variable_delay_unit_3.out VDPWR 1.34424f
C172 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VDPWR 0.706518f
C173 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 4.53e-19
C174 variable_delay_short_0.variable_delay_unit_2.out a_24240_17262# 0.505512f
C175 uo_out[4] uo_out[1] 2.26e-21
C176 uo_out[3] uo_out[2] 2.27264f
C177 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_2.out 0.235667f
C178 a_15680_14582# a_16500_14582# 0.004142f
C179 ui_in[5] a_25060_21092# 0.001909f
C180 a_12420_35540# uo_out[5] 0.013457f
C181 variable_delay_short_0.variable_delay_unit_3.out a_25060_18144# 0.070146f
C182 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VDPWR 0.706518f
C183 a_15322_7112# input_stage_0.fine_delay_unit_1.in 0.130264f
C184 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 1.99e-19
C185 a_13254_39726# uo_out[7] 0.188251f
C186 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 7.91e-21
C187 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.006183f
C188 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_4.out 0.235667f
C189 a_24240_20210# a_25060_20210# 0.004142f
C190 a_12420_32880# a_13254_32880# 0.003413f
C191 variable_delay_dummy_0.out input_stage_0.fine_delay_unit_1.in 0.024958f
C192 a_12310_28270# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.15e-21
C193 variable_delay_short_0.variable_delay_unit_2.in VDPWR 2.12807f
C194 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.120255f
C195 a_25060_18144# variable_delay_short_0.variable_delay_unit_2.in 7.65e-21
C196 a_23820_7082# ui_in[0] 0.003341f
C197 uio_in[5] a_16292_8080# 0.002587f
C198 a_12310_25988# a_12308_24168# 0.005984f
C199 ui_in[6] variable_delay_short_0.variable_delay_unit_2.out 0.224474f
C200 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_13254_35540# 0.012202f
C201 a_24240_15196# variable_delay_short_0.variable_delay_unit_1.in 7.65e-21
C202 variable_delay_short_0.out variable_delay_short_0.in 0.599483f
C203 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 5.04e-20
C204 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.014814f
C205 ui_in[1] variable_delay_short_0.variable_delay_unit_4.out 0.001119f
C206 ui_in[3] a_24240_21092# 0.001719f
C207 ui_in[4] ui_in[5] 3.94805f
C208 a_25060_20210# variable_delay_short_0.variable_delay_unit_3.in 8.82e-20
C209 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_13254_37444# 0.010872f
C210 variable_delay_short_0.variable_delay_unit_3.out a_24240_20210# 0.505512f
C211 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.start_buffer_0.start_delay 0.04313f
C212 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 6.08e-20
C213 a_12308_28732# a_12420_28694# 0.030083f
C214 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12308_28732# 2.36e-21
C215 ui_in[4] a_24240_26106# 0.00352f
C216 ui_in[4] a_24240_24040# 0.127858f
C217 tdc_0.diff_gen_0.delay_unit_2_6.in_1 VDPWR 4.42926f
C218 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_16500_11634# 2.39e-19
C219 input_stage_0.fine_delay_unit_0.in VDPWR 1.53841f
C220 a_25060_14314# ui_in[2] 3.98e-20
C221 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.754929f
C222 uo_out[7] tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.229856f
C223 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 a_12310_32834# 3.84e-19
C224 ui_in[6] uio_in[0] 9.78e-19
C225 a_9330_15214# VDPWR 1.15434f
C226 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.085059f
C227 uio_in[2] uio_in[5] 1.37e-20
C228 a_16500_12516# variable_delay_dummy_0.out 0.172055f
C229 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12310_30552# 0.196592f
C230 a_24240_17262# a_25060_17262# 0.004142f
C231 variable_delay_short_0.variable_delay_unit_3.in a_25060_17262# 0.054206f
C232 a_12310_32834# a_12308_31014# 0.005984f
C233 tdc_0.start_buffer_0.start_delay VDPWR 4.05162f
C234 a_25060_15196# VDPWR 0.001468f
C235 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_3.in 0.499092f
C236 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_13254_24130# 0.174293f
C237 a_10108_23452# a_12310_23706# 2.08e-21
C238 ui_in[7] variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 1.5e-19
C239 variable_delay_short_0.out a_16292_8344# 2.5e-19
C240 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.99e-19
C241 a_13254_30976# uo_out[3] 0.005542f
C242 uo_out[0] a_12310_23706# 0.098308f
C243 a_15680_15464# variable_delay_dummy_0.variable_delay_unit_1.in 7.65e-21
C244 a_24240_15196# variable_delay_short_0.variable_delay_unit_2.out 0.071074f
C245 a_12308_40142# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.100263f
C246 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.out 0.002141f
C247 a_16292_6966# uio_in[2] 0.024305f
C248 variable_delay_short_0.variable_delay_unit_4.out a_25060_23158# 0.222585f
C249 variable_delay_short_0.variable_delay_unit_5.in a_25060_23158# 0.054206f
C250 a_25060_24040# variable_delay_short_0.variable_delay_unit_4.in 7.65e-21
C251 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.6e-19
C252 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 VDPWR 5.07283f
C253 ui_in[5] ui_in[2] 7.13e-19
C254 uio_in[3] a_16292_8344# 0.025624f
C255 a_12308_26450# a_12310_28270# 0.005984f
C256 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12308_35578# 0.162625f
C257 a_23820_8460# variable_delay_short_0.out 0.00491f
C258 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.010157f
C259 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 VDPWR 5.07283f
C260 a_24240_17262# variable_delay_short_0.variable_delay_unit_2.in 8.82e-20
C261 input_stage_0.fine_delay_unit_0.in a_16292_8080# 1.39e-20
C262 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_2.in 0.087283f
C263 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.100263f
C264 tdc_0.diff_gen_0.delay_unit_2_6.in_2 tdc_0.diff_gen_0.delay_unit_2_5.in_2 0.04313f
C265 ui_in[6] a_25060_17262# 0.15982f
C266 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C267 ui_in[6] variable_delay_short_0.variable_delay_unit_3.out 0.043504f
C268 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_10108_32580# 0.09966f
C269 a_12308_33296# VDPWR 1.40782f
C270 uio_in[4] variable_delay_short_0.out 0.10432f
C271 ui_in[3] variable_delay_short_0.variable_delay_unit_4.in 0.02f
C272 a_16292_6702# input_stage_0.fine_delay_unit_1.in 7.4e-19
C273 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.006183f
C274 ui_in[7] a_25060_12248# 6.99e-20
C275 a_12420_35162# a_13254_35162# 0.003413f
C276 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14634# 0.00141f
C277 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.018644f
C278 a_13254_37822# VDPWR 6.18e-19
C279 uio_in[4] uio_in[3] 9.04698f
C280 a_15322_7112# uio_in[5] 0.007103f
C281 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.28924f
C282 a_24790_6672# ui_in[0] 0.022037f
C283 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_25060_20210# 2.39e-19
C284 input_stage_0.fine_delay_unit_0.in uio_in[2] 0.021403f
C285 ui_in[6] variable_delay_short_0.variable_delay_unit_2.in 0.50637f
C286 uio_in[5] variable_delay_dummy_0.out 0.126558f
C287 variable_delay_short_0.out input_stage_0.fine_delay_unit_1.in 0.008066f
C288 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.814958f
C289 uo_out[2] a_12308_28732# 0.014835f
C290 variable_delay_short_0.out variable_delay_short_0.variable_delay_unit_1.in 0.235655f
C291 a_9330_14634# VDPWR 1.15434f
C292 a_12420_35162# uo_out[5] 0.492009f
C293 uio_in[3] input_stage_0.fine_delay_unit_1.in 0.010396f
C294 uio_out[3] uio_out[2] 0.170937f
C295 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 3.26e-19
C296 ui_in[3] a_24240_11366# 0.001719f
C297 uio_out[5] uio_out[4] 0.170937f
C298 a_15322_7112# a_16292_6966# 0.019821f
C299 variable_delay_short_0.variable_delay_unit_4.out a_25060_21092# 0.070146f
C300 a_23820_7082# VDPWR 1.25441f
C301 a_24240_23158# variable_delay_short_0.variable_delay_unit_4.in 8.82e-20
C302 uio_out[7] uio_out[6] 0.170937f
C303 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.out 0.12029f
C304 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_5.in_2 0.401225f
C305 a_9330_15214# a_9330_15794# 0.001101f
C306 ui_in[7] ui_in[3] 0.014973f
C307 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.283838f
C308 a_24790_8050# variable_delay_short_0.out 6.1e-19
C309 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12310_35116# 0.164402f
C310 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_24240_12248# 0.029284f
C311 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_1.in 0.499092f
C312 a_24240_15196# variable_delay_short_0.variable_delay_unit_2.in 0.020173f
C313 a_12420_26034# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 1.47e-19
C314 a_24240_14314# VDPWR 1.6584f
C315 a_25060_15196# ui_in[6] 6.99e-20
C316 uio_in[1] VDPWR 6.39e-19
C317 a_24240_12248# variable_delay_short_0.in 7.65e-21
C318 ui_in[4] variable_delay_short_0.variable_delay_unit_5.in 0.607531f
C319 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_13254_28694# 0.174293f
C320 a_10108_28016# a_12310_28270# 2.08e-21
C321 ui_in[4] variable_delay_short_0.variable_delay_unit_4.out 0.227555f
C322 a_15322_7112# input_stage_0.fine_delay_unit_0.in 0.254311f
C323 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 VDPWR 3.23832f
C324 variable_delay_short_0.variable_delay_unit_5.forward a_25060_26106# 0.054206f
C325 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12310_23706# 0.196592f
C326 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12420_35540# 0.003607f
C327 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12310_25988# 0.196592f
C328 a_9330_15504# a_9330_15214# 0.083149f
C329 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 1.17e-19
C330 a_13254_40104# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.012202f
C331 uio_in[0] variable_delay_short_0.out 0.371181f
C332 input_stage_1.fine_delay_unit_1.in a_23820_7082# 0.130264f
C333 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 VDPWR 3.23832f
C334 a_12308_37860# a_13254_37822# 1.02e-19
C335 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12420_37822# 0.504416f
C336 ui_in[5] a_24240_18144# 6.99e-20
C337 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12310_23706# 0.014814f
C338 a_12310_30552# uo_out[3] 0.098308f
C339 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.in 0.499092f
C340 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.out 0.071795f
C341 a_9330_15214# tdc_0.diff_gen_0.delay_unit_2_2.in_2 5.93e-19
C342 a_12420_33258# VDPWR 0.497547f
C343 variable_delay_short_0.variable_delay_unit_4.in a_24240_21092# 0.020173f
C344 variable_delay_short_0.variable_delay_unit_5.forward ui_in[3] 0.007775f
C345 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 4.28924f
C346 a_16292_6702# uio_in[5] 9.94e-20
C347 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 uo_out[4] 0.20241f
C348 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VDPWR 0.706518f
C349 a_24240_15196# a_25060_15196# 0.011184f
C350 ui_in[5] variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 8.8e-19
C351 variable_delay_short_0.variable_delay_unit_5.in ui_in[2] 3.31e-20
C352 a_12308_31014# a_12420_30976# 0.030083f
C353 ui_in[2] variable_delay_short_0.variable_delay_unit_4.out 0.002549f
C354 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_1 0.001356f
C355 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_24240_24040# 0.029284f
C356 a_12420_26034# a_13254_26034# 0.003413f
C357 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_16500_14582# 2.39e-19
C358 variable_delay_short_0.variable_delay_unit_1.out uio_in[0] 0.043504f
C359 a_9330_14634# a_9330_15794# 2.78e-19
C360 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 0.231672f
C361 uio_in[5] variable_delay_short_0.out 0.082659f
C362 a_16292_6966# a_16292_6702# 0.556904f
C363 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq uo_out[4] 0.229249f
C364 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_10108_28016# 0.09966f
C365 uo_out[2] a_12420_28694# 0.013457f
C366 a_24790_6672# VDPWR 5.43e-20
C367 tdc_0.start_buffer_0.start_buff tdc_0.start_buffer_0.start_delay 1.12095f
C368 uo_out[3] VDPWR 0.587468f
C369 ui_in[4] a_25060_23158# 0.15982f
C370 ui_in[2] ui_in[1] 5.7665f
C371 uio_in[2] uio_in[1] 9.35827f
C372 uio_in[3] uio_in[5] 0.001464f
C373 ui_in[3] ui_in[0] 2.87e-19
C374 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 3.6e-19
C375 a_12310_37398# VDPWR 1.42789f
C376 a_24240_26988# ui_in[3] 0.001719f
C377 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 6.93e-19
C378 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 3.6e-19
C379 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 uo_out[3] 0.10528f
C380 variable_delay_dummy_0.variable_delay_unit_1.forward VDPWR 2.28565f
C381 a_13254_35162# uo_out[5] 0.188081f
C382 a_25060_14314# variable_delay_short_0.variable_delay_unit_1.in 8.82e-20
C383 variable_delay_short_0.variable_delay_unit_1.in a_24240_12248# 0.020173f
C384 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 5.04e-20
C385 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en VDPWR 2.77611f
C386 a_24790_8050# input_stage_1.fine_delay_unit_0.in 1.39e-20
C387 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VDPWR 0.706518f
C388 input_stage_0.fine_delay_unit_0.in a_16292_6702# 0.244525f
C389 ui_in[6] uio_in[1] 3.03e-19
C390 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_25060_18144# 0.15982f
C391 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_12308_28732# 5.04e-20
C392 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.010157f
C393 input_stage_1.fine_delay_unit_1.in a_24790_6672# 7.4e-19
C394 ui_in[2] a_25060_23158# 3.98e-20
C395 a_25284_5108# VDPWR 0.010256f
C396 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C397 uo_out[6] uo_out[4] 1.58e-19
C398 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[2] 6.97e-19
C399 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.in 0.235667f
C400 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.752988f
C401 variable_delay_dummy_0.variable_delay_unit_1.in a_16500_11634# 0.054206f
C402 ui_in[5] variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 7.3e-19
C403 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C404 a_9330_13764# VDPWR 1.15414f
C405 a_12420_37822# a_13254_37822# 0.003413f
C406 variable_delay_dummy_0.variable_delay_unit_1.forward a_15680_14582# 0.088132f
C407 uio_oe[4] uio_oe[3] 0.170937f
C408 a_15322_7112# uio_in[1] 0.003341f
C409 a_25060_12248# VDPWR 0.001468f
C410 tdc_0.start_buffer_0.start_delay variable_delay_short_0.out 6.15e-19
C411 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12310_28270# 0.014814f
C412 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_24240_26106# 0.11539f
C413 ui_in[4] a_25060_21092# 6.99e-20
C414 uio_in[1] variable_delay_dummy_0.out 0.001132f
C415 a_12308_24168# VDPWR 1.40782f
C416 uo_out[3] uo_out[1] 1.56e-19
C417 a_13254_35540# VDPWR 6.18e-19
C418 rst_n clk 0.031023f
C419 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12420_35162# 0.035356f
C420 tdc_0.diff_gen_0.delay_unit_2_3.in_2 VDPWR 3.06075f
C421 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.164402f
C422 a_12308_37860# a_12310_37398# 0.00595f
C423 a_12310_30552# a_12308_28732# 0.005984f
C424 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12420_37444# 0.013457f
C425 ui_in[5] variable_delay_short_0.variable_delay_unit_2.out 2.67e-19
C426 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 1.15e-21
C427 uio_in[4] variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.001173f
C428 uio_in[0] a_24240_12248# 0.124274f
C429 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_13254_33258# 0.012202f
C430 a_25060_26106# VDPWR 0.160518f
C431 a_25060_24040# VDPWR 0.001538f
C432 a_12420_32880# VDPWR 0.497771f
C433 a_13254_33258# uo_out[4] 0.005542f
C434 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.953579f
C435 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_24240_17262# 0.11539f
C436 a_25060_15196# variable_delay_short_0.variable_delay_unit_1.out 0.172055f
C437 ua[0] VDPWR 0.549361f
C438 variable_delay_short_0.variable_delay_unit_3.in variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.814958f
C439 uo_out[7] tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.105414f
C440 a_15680_11634# variable_delay_dummy_0.in 8.82e-20
C441 a_16500_15464# VDPWR 0.003377f
C442 ui_in[2] a_25060_21092# 3.98e-20
C443 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_13254_30976# 0.174293f
C444 a_12420_40104# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.003607f
C445 a_10108_30298# a_12310_30552# 2.08e-21
C446 uo_out[1] tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.229249f
C447 a_16786_5138# uio_in[5] 0.009499f
C448 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 uo_out[7] 1.53e-22
C449 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.out 0.12029f
C450 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 0.814958f
C451 a_24790_8314# ui_in[3] 0.024305f
C452 ui_in[3] VDPWR 0.206858f
C453 ui_in[5] uio_in[0] 3e-19
C454 a_25060_26988# variable_delay_short_0.variable_delay_unit_5.in 7.65e-21
C455 variable_delay_short_0.variable_delay_unit_5.out a_25060_26106# 0.222585f
C456 variable_delay_short_0.variable_delay_unit_5.out a_25060_24040# 0.070146f
C457 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 uo_out[2] 1.35e-20
C458 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.231672f
C459 ui_in[3] a_25060_18144# 0.002391f
C460 uo_out[2] a_12420_28316# 0.492009f
C461 a_12308_28732# VDPWR 1.40782f
C462 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_12308_40142# 0.197073f
C463 ui_in[6] variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 1.09842f
C464 a_9330_14634# variable_delay_short_0.out 2.11e-19
C465 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 3.26e-19
C466 ui_in[5] a_25060_20210# 0.15982f
C467 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 4.53e-19
C468 tdc_0.diff_gen_0.delay_unit_2_3.in_1 VDPWR 4.44087f
C469 a_13254_26412# VDPWR 6.18e-19
C470 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.010157f
C471 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq uo_out[6] 0.229249f
C472 variable_delay_short_0.variable_delay_unit_5.out ui_in[3] 0.040959f
C473 uo_out[0] uio_in[5] 1.28234f
C474 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12308_37860# 0.197073f
C475 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12308_28732# 3.26e-19
C476 ui_in[4] ui_in[2] 7.13e-19
C477 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 1.17e-19
C478 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.6e-19
C479 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14924# 6.93e-19
C480 uo_out[1] a_12308_24168# 6.49e-20
C481 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_12308_33296# 0.162625f
C482 a_16292_6702# uio_in[1] 0.022338f
C483 a_25060_14314# variable_delay_short_0.variable_delay_unit_2.in 0.054206f
C484 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 VDPWR 3.23832f
C485 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.871529f
C486 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.002365f
C487 a_12420_37444# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 1.47e-19
C488 a_24240_23158# VDPWR 1.6584f
C489 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_16500_12516# 0.15982f
C490 ui_in[5] variable_delay_short_0.variable_delay_unit_3.out 0.22469f
C491 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_10108_30298# 0.09966f
C492 ui_in[3] a_24240_20210# 0.001719f
C493 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.59e-20
C494 input_stage_1.fine_delay_unit_1.in ui_in[3] 0.020481f
C495 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 0.100263f
C496 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_12420_28316# 1.47e-19
C497 a_9330_14924# VDPWR 1.1544f
C498 variable_delay_dummy_0.variable_delay_unit_1.out uio_in[4] 4.58e-20
C499 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 a_12308_31014# 5.04e-20
C500 uio_in[1] variable_delay_short_0.out 0.030581f
C501 a_12420_24130# VDPWR 0.497547f
C502 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 9.61e-20
C503 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.002365f
C504 tdc_0.diff_gen_0.delay_unit_2_3.in_2 a_9330_15794# 0.00105f
C505 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_25060_23158# 2.39e-19
C506 uio_in[3] uio_in[1] 0.001793f
C507 ui_in[3] a_24240_17262# 0.001719f
C508 ui_in[3] variable_delay_short_0.variable_delay_unit_3.in 0.02f
C509 uio_in[5] uio_in[6] 0.073214f
C510 input_stage_0.nand_gate_0.out uio_in[5] 0.283562f
C511 a_15680_11634# VDPWR 1.70112f
C512 a_12420_23752# a_13254_23752# 0.003413f
C513 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.out 0.002141f
C514 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.in 0.09141f
C515 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_10108_25734# 1.06381f
C516 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 6.93e-19
C517 variable_delay_short_0.variable_delay_unit_1.out a_24240_14314# 0.505512f
C518 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_13254_35162# 0.010872f
C519 a_12310_35116# VDPWR 1.42789f
C520 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_2 0.04313f
C521 uo_out[6] tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 1.35e-20
C522 ui_in[2] a_25060_11366# 3.98e-20
C523 a_16292_6966# input_stage_0.nand_gate_0.out 4.47e-20
C524 uo_out[1] a_13254_26412# 0.005542f
C525 a_23820_7082# a_24790_6936# 0.019821f
C526 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.6e-19
C527 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_13254_37444# 0.005542f
C528 ui_in[6] ui_in[3] 0.014973f
C529 uio_in[5] variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.026424f
C530 a_24240_21092# VDPWR 1.6584f
C531 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_12310_32834# 0.164402f
C532 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_13254_28694# 0.012202f
C533 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 uo_out[2] 3.69e-19
C534 a_12310_32834# uo_out[4] 0.098308f
C535 a_13254_32880# VDPWR 6.18e-19
C536 a_12420_28694# VDPWR 0.497547f
C537 tdc_0.start_buffer_0.start_buff a_9330_13764# 5.99e-19
C538 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.04313f
C539 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C540 a_9330_14634# a_9330_14344# 0.083149f
C541 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 uo_out[5] 0.20241f
C542 a_10108_25734# a_12310_25988# 2.08e-21
C543 uio_out[2] uio_out[1] 0.170937f
C544 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 1.17e-19
C545 variable_delay_dummy_0.variable_delay_unit_1.out a_16500_12516# 0.070146f
C546 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12310_30552# 0.014814f
C547 a_13254_37822# uo_out[6] 0.005542f
C548 a_12420_39726# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.035356f
C549 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 5.04e-20
C550 uio_out[6] uio_out[5] 0.170937f
C551 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12420_37822# 0.033952f
C552 a_24790_8050# ui_in[1] 7.45e-19
C553 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 4.53e-19
C554 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 a_12308_24168# 5.04e-20
C555 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_12420_33258# 0.003607f
C556 a_23820_7082# input_stage_1.fine_delay_unit_0.in 0.254311f
C557 uo_out[2] a_13254_28316# 0.188081f
C558 input_stage_0.fine_delay_unit_0.in input_stage_0.nand_gate_0.out 0.062023f
C559 ui_in[1] variable_delay_short_0.variable_delay_unit_2.out 0.001119f
C560 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.59e-20
C561 tdc_0.diff_gen_0.delay_unit_2_4.in_2 tdc_0.diff_gen_0.delay_unit_2_3.in_1 0.311186f
C562 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_2 0.401225f
C563 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.100263f
C564 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.138497f
C565 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C566 a_24240_15196# ui_in[3] 0.001719f
C567 a_9330_14924# a_9330_15794# 4.98e-19
C568 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 uo_out[4] 1.35e-20
C569 uio_in[4] a_16500_11634# 6.61e-20
C570 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_1.in 0.09141f
C571 a_12310_25988# VDPWR 1.42789f
C572 ui_in[3] variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 0.014554f
C573 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.953579f
C574 variable_delay_dummy_0.variable_delay_unit_1.out a_16500_14582# 0.222585f
C575 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12420_33258# 0.504416f
C576 a_12308_33296# a_13254_33258# 1.02e-19
C577 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_12308_31014# 3.26e-19
C578 ui_in[4] variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 1.11761f
C579 a_12308_31014# uo_out[4] 6.49e-20
C580 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VDPWR 0.706518f
C581 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12308_28732# 0.162625f
C582 ui_in[4] a_25060_26988# 8.92e-19
C583 tdc_0.vernier_delay_line_0.start_neg VDPWR 3.22778f
C584 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.401225f
C585 tdc_0.diff_gen_0.delay_unit_2_3.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.311186f
C586 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_10108_39426# 1.06381f
C587 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.forward 0.794183f
C588 a_24240_26988# variable_delay_short_0.variable_delay_unit_5.forward 0.016896f
C589 ui_in[2] variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 6.97e-19
C590 variable_delay_short_0.variable_delay_unit_4.in VDPWR 2.12807f
C591 a_12308_35578# a_12310_37398# 0.005984f
C592 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.231672f
C593 a_24240_21092# variable_delay_short_0.variable_delay_unit_3.in 7.65e-21
C594 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_10108_37144# 1.06381f
C595 variable_delay_dummy_0.variable_delay_unit_1.out uio_in[5] 0.016377f
C596 a_9330_13764# variable_delay_short_0.out 0.076613f
C597 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.out 0.071795f
C598 ui_in[2] variable_delay_short_0.in 1.86e-20
C599 a_12420_28316# a_13254_28316# 0.003413f
C600 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 a_12420_30598# 1.47e-19
C601 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 4.53e-19
C602 a_23820_7082# input_stage_1.nand_gate_0.out 3.78e-19
C603 variable_delay_short_0.out a_25060_12248# 0.172055f
C604 a_24790_6936# a_24790_6672# 0.556904f
C605 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.002141f
C606 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.out 0.085059f
C607 a_12420_23752# VDPWR 0.497771f
C608 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.018644f
C609 a_24240_14314# a_25060_14314# 0.004142f
C610 uo_out[1] tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.20241f
C611 a_9330_14054# a_9330_13764# 0.083149f
C612 uo_out[2] VDPWR 0.587468f
C613 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_3.in_1 0.756572f
C614 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.231672f
C615 uo_out[6] tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 3.69e-19
C616 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_25060_11366# 2.39e-19
C617 ui_in[2] variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 6.97e-19
C618 a_12420_37444# a_12310_37398# 0.030392f
C619 a_25060_26988# ui_in[2] 3.98e-20
C620 ui_in[1] variable_delay_short_0.variable_delay_unit_3.out 0.001119f
C621 a_25060_11366# variable_delay_short_0.in 8.82e-20
C622 a_24240_11366# VDPWR 1.6584f
C623 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 uo_out[2] 6.28e-22
C624 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en uio_in[0] 1.5e-19
C625 variable_delay_dummy_0.out a_15680_11634# 0.505512f
C626 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.003768f
C627 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.756572f
C628 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 a_10108_32580# 0.007929f
C629 ui_in[5] uio_in[1] 1.46e-19
C630 variable_delay_short_0.variable_delay_unit_4.in a_24240_20210# 0.088132f
C631 tdc_0.start_buffer_0.start_delay a_7140_10670# 7.1e-20
C632 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_12308_24168# 0.197073f
C633 variable_delay_short_0.variable_delay_unit_1.out a_25060_12248# 0.070146f
C634 uo_out[1] a_12310_25988# 0.098308f
C635 input_stage_1.fine_delay_unit_0.in a_24790_6672# 0.244525f
C636 uio_in[4] variable_delay_dummy_0.variable_delay_unit_1.in 4.58e-20
C637 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 3.26e-19
C638 ui_in[7] VDPWR 1.41097f
C639 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.626611f
C640 a_23820_8460# ui_in[2] 0.003402f
C641 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_12308_24168# 3.26e-19
C642 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 VDPWR 5.07283f
C643 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12310_28270# 0.164402f
C644 ui_in[3] variable_delay_short_0.out 0.06888f
C645 a_12420_28316# VDPWR 0.497771f
C646 ui_in[4] variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en 0.025512f
C647 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.953579f
C648 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_3.in 0.087283f
C649 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 uo_out[5] 1.53e-22
C650 a_12308_35578# a_13254_35540# 1.02e-19
C651 uo_out[6] uo_out[3] 2.26e-21
C652 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12420_35540# 0.504416f
C653 uo_out[5] uo_out[4] 1.5647f
C654 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_16500_15464# 0.15982f
C655 a_12310_37398# uo_out[6] 0.098308f
C656 a_13254_39726# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.010872f
C657 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_24240_21092# 0.029284f
C658 a_12420_35162# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 1.47e-19
C659 input_stage_0.nand_gate_0.out uio_in[1] 1.7e-19
C660 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 6.93e-19
C661 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12420_37444# 0.003664f
C662 a_12420_33258# a_13254_33258# 0.003413f
C663 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 a_12420_23752# 1.47e-19
C664 a_13254_30976# VDPWR 6.18e-19
C665 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.100263f
C666 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_12420_32880# 0.035356f
C667 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12420_28694# 0.003607f
C668 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 3.6e-19
C669 uo_out[2] uo_out[1] 2.62662f
C670 uo_out[3] uo_out[0] 2.26e-21
C671 uio_in[5] a_16500_11634# 0.002787f
C672 ui_in[6] variable_delay_short_0.variable_delay_unit_4.in 0.001632f
C673 variable_delay_short_0.variable_delay_unit_1.out ui_in[3] 0.040959f
C674 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.in 0.814958f
C675 a_24790_6672# input_stage_1.nand_gate_0.out 5.26e-20
C676 variable_delay_short_0.variable_delay_unit_5.forward VDPWR 2.28561f
C677 ui_in[2] variable_delay_short_0.variable_delay_unit_1.in 3.31e-20
C678 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_13254_30976# 0.012202f
C679 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.45e-19
C680 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en ui_in[2] 6.97e-19
C681 uio_oe[3] uio_oe[2] 0.170937f
C682 a_12308_33296# a_12310_32834# 0.00595f
C683 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12420_32880# 0.013457f
C684 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.in 0.091118f
C685 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.006183f
C686 a_9330_14924# variable_delay_short_0.out 8.85e-20
C687 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.132512f
C688 ui_in[7] uio_in[2] 2.48e-19
C689 uo_out[6] tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 6.28e-22
C690 clk ena 0.031023f
C691 ui_in[4] uio_in[0] 1.15e-19
C692 variable_delay_dummy_0.in a_15322_8490# 0.123564f
C693 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.forward 0.234428f
C694 a_13254_26412# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.012202f
C695 ui_in[7] variable_delay_short_0.variable_delay_unit_3.in 3.37e-20
C696 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 2.59e-20
C697 variable_delay_short_0.variable_delay_unit_1.in a_25060_11366# 0.054206f
C698 a_9330_15214# tdc_0.diff_gen_0.delay_unit_2_1.in_1 5.9e-19
C699 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 uo_out[6] 0.10528f
C700 a_24790_8050# ui_in[2] 0.023539f
C701 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.132512f
C702 a_25060_21092# variable_delay_short_0.variable_delay_unit_3.out 0.172055f
C703 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.752988f
C704 tdc_0.start_buffer_0.start_delay tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.401491f
C705 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.59e-20
C706 ui_in[0] VDPWR 6.58e-19
C707 ui_in[5] variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 9.38e-20
C708 a_13254_23752# VDPWR 6.18e-19
C709 ui_in[2] variable_delay_short_0.variable_delay_unit_2.out 0.002549f
C710 a_24240_26988# VDPWR 1.78268f
C711 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 9.61e-20
C712 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.010157f
C713 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 0.814958f
C714 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_12420_24130# 0.033952f
C715 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_25060_15196# 0.15982f
C716 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.2373f
C717 a_15680_15464# variable_delay_dummy_0.variable_delay_unit_1.forward 0.016896f
C718 a_16500_14582# variable_delay_dummy_0.variable_delay_unit_1.in 8.82e-20
C719 input_stage_1.nand_gate_0.out a_25284_5108# 0.355469f
C720 a_24240_12248# a_25060_12248# 0.011184f
C721 a_13254_40104# VDPWR 6.18e-19
C722 ui_in[6] ui_in[7] 7.62803f
C723 a_12310_37398# a_13254_37444# 1.02e-19
C724 input_stage_1.fine_delay_unit_0.in ua[0] 5.53e-19
C725 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12308_31014# 0.162625f
C726 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.019727f
C727 variable_delay_dummy_0.in VDPWR 1.61964f
C728 a_24240_26988# variable_delay_short_0.variable_delay_unit_5.out 0.493816f
C729 a_15680_12516# variable_delay_dummy_0.in 7.65e-21
C730 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 VDPWR 3.23832f
C731 uo_out[0] a_12308_24168# 0.014835f
C732 uio_in[0] ui_in[2] 7.13e-19
C733 ui_in[4] variable_delay_short_0.variable_delay_unit_3.out 2.67e-19
C734 a_16786_5138# ua[0] 0.009499f
C735 uo_out[2] tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.20241f
C736 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 1.24e-19
C737 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 6.93e-19
C738 a_23820_8460# variable_delay_short_0.in 0.121301f
C739 a_23820_7082# ui_in[1] 0.010812f
C740 a_12420_35540# a_13254_35540# 0.003413f
C741 uio_in[5] variable_delay_dummy_0.variable_delay_unit_1.in 0.019965f
C742 a_12420_30598# a_13254_30598# 0.003413f
C743 ui_in[2] a_25060_20210# 3.98e-20
C744 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.018644f
C745 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12420_26412# 0.504416f
C746 a_12308_26450# a_13254_26412# 1.02e-19
C747 uio_in[0] a_25060_11366# 0.15982f
C748 a_13254_28316# VDPWR 6.18e-19
C749 a_12310_35116# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.45e-19
C750 a_24240_15196# ui_in[7] 0.124274f
C751 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 4.53e-19
C752 a_12308_35578# a_12310_35116# 0.00595f
C753 a_25060_14314# ui_in[3] 0.002391f
C754 variable_delay_dummy_0.in a_16292_8080# 3.44e-20
C755 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12420_35162# 0.013457f
C756 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 6.79e-20
C757 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 7.91e-21
C758 ui_in[3] a_24240_12248# 0.001719f
C759 ui_in[6] variable_delay_short_0.variable_delay_unit_5.forward 0.001598f
C760 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.814958f
C761 ui_in[2] a_25060_17262# 3.98e-20
C762 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.499806f
C763 input_stage_1.nand_gate_0.out ua[0] 0.050326f
C764 a_13254_40104# uo_out[7] 0.005712f
C765 ui_in[2] variable_delay_short_0.variable_delay_unit_3.out 0.002549f
C766 a_24240_26106# a_25060_26106# 0.004142f
C767 a_24240_24040# a_25060_24040# 0.011184f
C768 a_15322_8490# VDPWR 1.25073f
C769 a_12310_30552# VDPWR 1.42789f
C770 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 4.53e-19
C771 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 4.28924f
C772 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.499806f
C773 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_13254_32880# 0.010872f
C774 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_12420_28316# 0.035356f
C775 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.in 0.08442f
C776 a_12310_35116# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 6.08e-20
C777 ui_in[5] ui_in[3] 0.014973f
C778 tdc_0.diff_gen_0.delay_unit_2_1.in_2 VDPWR 3.06163f
C779 uio_in[2] variable_delay_dummy_0.in 1.05e-20
C780 uio_in[4] a_16292_8344# 0.024305f
C781 a_15680_15464# a_16500_15464# 0.011184f
C782 ui_in[2] variable_delay_short_0.variable_delay_unit_2.in 3.31e-20
C783 a_12420_40104# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.504416f
C784 a_13254_40104# a_12308_40142# 1.02e-19
C785 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 uo_out[5] 1.35e-20
C786 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12310_30552# 0.164402f
C787 a_24240_26106# ui_in[3] 0.001719f
C788 ui_in[3] a_24240_24040# 0.001719f
C789 a_12310_25988# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 1.15e-21
C790 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.283838f
C791 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 0.002365f
C792 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_13254_32880# 0.005542f
C793 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_25060_26988# 0.15982f
C794 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 2.59e-20
C795 a_12308_33296# uo_out[5] 6.49e-20
C796 input_stage_0.nand_gate_0.out ua[0] 0.050326f
C797 tdc_0.vernier_delay_line_0.start_neg tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.007279f
C798 a_24790_8050# variable_delay_short_0.in 3.44e-20
C799 a_15322_8490# a_16292_8080# 0.53267f
C800 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.747722f
C801 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_24240_14314# 0.11539f
C802 a_12310_25988# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.164402f
C803 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 6.79e-20
C804 input_stage_0.fine_delay_unit_1.in a_16292_8344# 0.028846f
C805 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12308_35578# 0.197073f
C806 a_15680_12516# VDPWR 1.78275f
C807 a_25060_18144# VDPWR 0.001468f
C808 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12420_30976# 0.003607f
C809 a_24240_18144# variable_delay_short_0.variable_delay_unit_2.out 0.493816f
C810 a_24790_6672# ui_in[1] 0.00799f
C811 variable_delay_short_0.out a_24240_11366# 0.505512f
C812 uio_in[0] variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 1.09349f
C813 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C814 uo_out[0] a_12420_24130# 0.013457f
C815 variable_delay_short_0.variable_delay_unit_5.out VDPWR 1.5668f
C816 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.018644f
C817 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_12420_23752# 0.003664f
C818 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.variable_delay_unit_1.forward 0.234428f
C819 uio_in[4] input_stage_0.fine_delay_unit_1.in 0.020481f
C820 uio_out[1] uio_out[0] 0.170937f
C821 a_25060_15196# ui_in[2] 3.98e-20
C822 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12308_26450# 0.162625f
C823 uio_in[0] variable_delay_short_0.in 0.26219f
C824 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12308_24168# 0.162625f
C825 a_12310_39680# VDPWR 1.42789f
C826 a_15680_14582# VDPWR 1.70112f
C827 ui_in[7] variable_delay_short_0.out 2.67e-19
C828 a_12420_26412# a_13254_26412# 0.003413f
C829 a_12308_24168# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.100263f
C830 a_12308_31014# uo_out[3] 0.014835f
C831 variable_delay_dummy_0.out variable_delay_dummy_0.in 0.728538f
C832 uo_out[2] tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.53e-22
C833 a_24240_20210# VDPWR 1.6584f
C834 a_23820_8460# a_24790_8050# 0.53267f
C835 input_stage_1.fine_delay_unit_1.in a_24790_8314# 0.028846f
C836 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.006183f
C837 input_stage_1.fine_delay_unit_1.in VDPWR 1.33479f
C838 ui_in[7] uio_in[3] 1.26e-19
C839 uo_out[7] VDPWR 0.587468f
C840 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.2373f
C841 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.006183f
C842 a_12308_26450# a_12310_25988# 0.00595f
C843 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12420_26034# 0.013457f
C844 uio_in[2] VDPWR 0.005628f
C845 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.2373f
C846 uio_in[4] a_16500_12516# 6.61e-20
C847 a_24240_17262# VDPWR 1.6584f
C848 a_12420_39726# a_13254_39726# 0.003413f
C849 variable_delay_short_0.variable_delay_unit_3.in VDPWR 2.12807f
C850 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 VDPWR 5.20504f
C851 a_12308_40142# VDPWR 1.40742f
C852 variable_delay_short_0.variable_delay_unit_1.out ui_in[7] 0.224474f
C853 uo_out[1] VDPWR 0.587468f
C854 ui_in[5] a_24240_21092# 0.124669f
C855 a_23820_8460# uio_in[0] 1.26e-19
C856 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13254_35162# 0.005542f
C857 variable_delay_short_0.variable_delay_unit_3.out a_24240_18144# 0.071074f
C858 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 0.031607f
C859 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 uo_out[6] 1.53e-22
C860 a_12308_37860# VDPWR 1.40782f
C861 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.in 7.91e-21
C862 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 uo_out[5] 3.69e-19
C863 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 2.59e-20
C864 a_12310_39680# uo_out[7] 0.098487f
C865 a_15322_7112# a_15322_8490# 0.001571f
C866 a_25060_24040# variable_delay_short_0.variable_delay_unit_4.out 0.172055f
C867 a_25060_26106# variable_delay_short_0.variable_delay_unit_5.in 8.82e-20
C868 a_12420_32880# a_12310_32834# 0.030392f
C869 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.003768f
C870 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.out 0.002141f
C871 variable_delay_dummy_0.out a_15322_8490# 0.011089f
C872 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.499806f
C873 a_9330_15794# VDPWR 1.86061f
C874 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_13254_28316# 0.010872f
C875 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.002365f
C876 tdc_0.diff_gen_0.delay_unit_2_5.in_2 VDPWR 3.06042f
C877 a_24240_18144# variable_delay_short_0.variable_delay_unit_2.in 7.65e-21
C878 ui_in[6] VDPWR 1.41131f
C879 uio_in[5] a_16292_8344# 0.001923f
C880 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq uo_out[5] 0.229249f
C881 ui_in[6] a_25060_18144# 0.001909f
C882 uio_in[2] a_16292_8080# 0.001529f
C883 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12420_35540# 0.033952f
C884 a_16500_15464# variable_delay_dummy_0.variable_delay_unit_1.out 0.172055f
C885 uo_out[2] a_12308_26450# 6.49e-20
C886 a_12420_39726# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.013457f
C887 a_12310_39680# a_12308_40142# 0.00595f
C888 variable_delay_short_0.variable_delay_unit_5.in ui_in[3] 0.02f
C889 ui_in[3] variable_delay_short_0.variable_delay_unit_4.out 0.040959f
C890 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12310_37398# 0.196592f
C891 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 3.45e-19
C892 a_24240_20210# variable_delay_short_0.variable_delay_unit_3.in 8.82e-20
C893 a_12310_39680# a_12308_37860# 0.005984f
C894 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_15680_11634# 0.11539f
C895 uio_in[0] variable_delay_short_0.variable_delay_unit_1.in 0.574722f
C896 tdc_0.diff_gen_0.delay_unit_2_4.in_2 VDPWR 3.06175f
C897 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.04313f
C898 a_15322_7112# VDPWR 1.25441f
C899 uo_out[7] a_12308_40142# 0.01561f
C900 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 a_12420_32880# 1.47e-19
C901 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 uo_out[4] 0.10528f
C902 a_9330_15504# VDPWR 1.1544f
C903 uo_out[5] uo_out[3] 1.56e-19
C904 variable_delay_dummy_0.out VDPWR 1.79065f
C905 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12420_26412# 0.003607f
C906 uio_in[4] uio_in[5] 7.75329f
C907 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12420_24130# 0.003607f
C908 ui_in[3] ui_in[1] 0.018155f
C909 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 8.54e-19
C910 a_15680_12516# variable_delay_dummy_0.out 0.493816f
C911 a_12308_37860# uo_out[7] 6.49e-20
C912 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12420_30598# 0.035356f
C913 variable_delay_short_0.variable_delay_unit_3.in a_24240_17262# 0.088132f
C914 a_24240_15196# VDPWR 1.6584f
C915 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.start_buffer_0.start_buff 0.311237f
C916 a_12308_24168# a_13254_24130# 1.02e-19
C917 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12420_24130# 0.504416f
C918 ui_in[5] variable_delay_short_0.variable_delay_unit_4.in 0.586739f
C919 tdc_0.diff_gen_0.delay_unit_2_2.in_2 VDPWR 3.0616f
C920 a_12308_28732# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.100263f
C921 a_12420_30976# uo_out[3] 0.013457f
C922 variable_delay_short_0.out variable_delay_dummy_0.in 0.100566f
C923 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en VDPWR 2.77611f
C924 uo_out[0] a_12420_23752# 0.492009f
C925 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C926 uo_out[7] uio_out[0] 0.170937f
C927 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 a_12310_32834# 4.55e-19
C928 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 4.28924f
C929 uo_out[2] uo_out[0] 1.56e-19
C930 variable_delay_short_0.variable_delay_unit_4.out a_24240_23158# 0.505512f
C931 variable_delay_short_0.variable_delay_unit_5.in a_24240_23158# 0.088132f
C932 a_24240_24040# variable_delay_short_0.variable_delay_unit_4.in 7.65e-21
C933 uio_in[5] input_stage_0.fine_delay_unit_1.in 0.011377f
C934 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_10108_34862# 1.06381f
C935 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.010157f
C936 uio_in[3] variable_delay_dummy_0.in 5.31e-20
C937 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.747722f
C938 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 6.79e-20
C939 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.499806f
C940 tdc_0.start_buffer_0.start_buff VDPWR 7.34803f
C941 ui_in[6] uio_in[2] 1.69e-19
C942 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.747722f
C943 ui_in[6] a_24240_17262# 0.042718f
C944 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 4.28924f
C945 variable_delay_dummy_0.out a_16292_8080# 6.96e-19
C946 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 6.79e-20
C947 ui_in[6] variable_delay_short_0.variable_delay_unit_3.in 0.580889f
C948 tdc_0.diff_gen_0.delay_unit_2_4.in_1 VDPWR 4.44109f
C949 ui_in[3] a_25060_23158# 0.002391f
C950 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.401225f
C951 a_25060_14314# ui_in[7] 0.15982f
C952 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 VDPWR 3.23844f
C953 a_16292_6966# input_stage_0.fine_delay_unit_1.in 5.97e-19
C954 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12308_33296# 7.19e-22
C955 a_12420_35162# a_12310_35116# 0.030392f
C956 ui_in[7] a_24240_12248# 6.99e-20
C957 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[3] 0.014554f
C958 a_12420_37822# VDPWR 0.497547f
C959 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 3.6e-19
C960 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.953579f
C961 variable_delay_short_0.variable_delay_unit_1.in variable_delay_short_0.variable_delay_unit_2.in 0.087283f
C962 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 uo_out[5] 6.28e-22
C963 tdc_0.diff_gen_0.delay_unit_2_3.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.001356f
C964 a_24790_6936# ui_in[0] 0.022567f
C965 uio_oe[2] uio_oe[1] 0.170937f
C966 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_24240_20210# 0.11539f
C967 a_15322_7112# uio_in[2] 0.010812f
C968 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 9.61e-20
C969 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_13254_26034# 0.005542f
C970 variable_delay_dummy_0.variable_delay_unit_1.forward variable_delay_dummy_0.variable_delay_unit_1.in 0.087283f
C971 uio_in[5] a_16500_12516# 0.002787f
C972 variable_delay_short_0.out a_15322_8490# 7.6e-19
C973 tdc_0.diff_gen_0.delay_unit_2_2.in_1 VDPWR 4.44107f
C974 uio_in[2] variable_delay_dummy_0.out 0.001744f
C975 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.2373f
C976 ui_in[5] ui_in[7] 0.00231f
C977 variable_delay_short_0.variable_delay_unit_2.out a_25060_17262# 0.222585f
C978 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.out 0.071795f
C979 a_13254_35540# uo_out[5] 0.005542f
C980 uio_in[3] a_15322_8490# 0.003646f
C981 variable_delay_short_0.variable_delay_unit_4.out a_24240_21092# 0.071074f
C982 input_stage_0.fine_delay_unit_0.in input_stage_0.fine_delay_unit_1.in 0.029975f
C983 a_24240_23158# a_25060_23158# 0.004142f
C984 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.in 0.09141f
C985 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_2 0.04313f
C986 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14054# 8.73e-19
C987 a_12310_32834# a_13254_32880# 1.02e-19
C988 a_12310_25988# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 3.45e-19
C989 a_9330_14924# tdc_0.diff_gen_0.delay_unit_2_1.in_1 2.18e-19
C990 a_9330_15504# a_9330_15794# 0.087529f
C991 ui_in[2] variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 6.97e-19
C992 variable_delay_short_0.variable_delay_unit_2.out variable_delay_short_0.variable_delay_unit_2.in 0.499092f
C993 input_stage_1.fine_delay_unit_0.in ui_in[0] 0.009426f
C994 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 uo_out[3] 1.35e-20
C995 a_12310_25988# tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 6.08e-20
C996 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12420_35162# 0.003664f
C997 a_24790_8314# variable_delay_short_0.out 4.38e-19
C998 variable_delay_short_0.out VDPWR 1.72578f
C999 a_25060_15196# variable_delay_short_0.variable_delay_unit_1.in 7.65e-21
C1000 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 1.24e-19
C1001 ui_in[3] a_25060_21092# 0.002391f
C1002 a_13254_39726# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.005542f
C1003 tdc_0.diff_gen_0.delay_unit_2_2.in_2 a_9330_15794# 0.001232f
C1004 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.192064f
C1005 a_24240_15196# ui_in[6] 6.99e-20
C1006 a_9330_14054# VDPWR 1.1544f
C1007 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.953579f
C1008 a_12420_24130# a_13254_24130# 0.003413f
C1009 variable_delay_short_0.variable_delay_unit_3.out a_25060_20210# 0.222585f
C1010 ui_in[6] variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 4.42e-19
C1011 uio_in[3] VDPWR 0.001248f
C1012 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_10108_28016# 0.192064f
C1013 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.09966f
C1014 ui_in[5] variable_delay_short_0.variable_delay_unit_5.forward 0.003308f
C1015 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 2.59e-20
C1016 a_12308_28732# a_13254_28694# 1.02e-19
C1017 ui_in[4] a_25060_24040# 0.001909f
C1018 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12420_28694# 0.504416f
C1019 uio_in[0] variable_delay_short_0.variable_delay_unit_2.in 3.37e-20
C1020 tdc_0.vernier_delay_line_0.start_pos tdc_0.diff_gen_0.delay_unit_2_6.in_2 0.400636f
C1021 variable_delay_short_0.variable_delay_unit_5.forward a_24240_26106# 0.088132f
C1022 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en VDPWR 3.86972f
C1023 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 1.17e-19
C1024 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12420_26034# 0.035356f
C1025 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_12420_23752# 0.035356f
C1026 ui_in[2] a_25060_12248# 3.98e-20
C1027 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43941f
C1028 a_23820_8460# a_23820_7082# 0.001571f
C1029 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_13254_30598# 0.010872f
C1030 a_12420_40104# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.033952f
C1031 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.2373f
C1032 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 6.08e-20
C1033 a_12308_37860# a_12420_37822# 0.030083f
C1034 ui_in[4] ui_in[3] 2.58276f
C1035 variable_delay_short_0.variable_delay_unit_1.out VDPWR 1.34424f
C1036 tdc_0.diff_gen_0.delay_unit_2_5.in_2 tdc_0.diff_gen_0.delay_unit_2_4.in_1 0.311186f
C1037 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_12420_23752# 0.013457f
C1038 a_12308_24168# a_12310_23706# 0.00595f
C1039 variable_delay_short_0.out a_16292_8080# 3.3e-19
C1040 a_12420_30598# uo_out[3] 0.492009f
C1041 uo_out[0] a_13254_23752# 0.188081f
C1042 a_16500_15464# variable_delay_dummy_0.variable_delay_unit_1.in 7.65e-21
C1043 a_25060_15196# variable_delay_short_0.variable_delay_unit_2.out 0.070146f
C1044 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 VDPWR 2.43248f
C1045 a_9330_15504# tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.001226f
C1046 input_stage_1.nand_gate_0.out ui_in[0] 1.7e-19
C1047 a_16292_6966# uio_in[5] 2.26e-20
C1048 a_16292_6702# uio_in[2] 0.00799f
C1049 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_4.in 0.499092f
C1050 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C1051 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_4.in 0.087283f
C1052 a_12308_35578# VDPWR 1.40782f
C1053 a_15680_11634# a_16500_11634# 0.004142f
C1054 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.132512f
C1055 input_stage_1.fine_delay_unit_1.in variable_delay_short_0.out 0.024792f
C1056 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_12310_28270# 6.08e-20
C1057 uio_in[3] a_16292_8080# 0.023966f
C1058 ui_in[5] a_24240_26988# 2.89e-20
C1059 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 6.93e-19
C1060 a_25060_26106# ui_in[2] 3.98e-20
C1061 ui_in[2] a_25060_24040# 3.98e-20
C1062 a_25060_17262# variable_delay_short_0.variable_delay_unit_2.in 8.82e-20
C1063 tdc_0.diff_gen_0.delay_unit_2_2.in_1 a_9330_15794# 4.02e-19
C1064 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.003768f
C1065 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_4.in_2 0.667766f
C1066 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_15680_14582# 0.11539f
C1067 tdc_0.start_buffer_0.start_buff variable_delay_dummy_0.out 5.26e-19
C1068 a_12420_26034# a_12310_25988# 0.030392f
C1069 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 6.79e-20
C1070 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.747722f
C1071 uio_in[2] variable_delay_short_0.out 0.022033f
C1072 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_12308_33296# 0.197073f
C1073 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VDPWR 0.706518f
C1074 a_12308_33296# uo_out[4] 0.014835f
C1075 uo_out[3] tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.53e-22
C1076 tdc_0.vernier_delay_line_0.start_pos tdc_0.diff_gen_0.delay_unit_2_6.in_1 0.728719f
C1077 a_12310_35116# a_13254_35162# 1.02e-19
C1078 tdc_0.diff_gen_0.delay_unit_2_1.in_2 a_9330_14344# 0.001157f
C1079 ui_in[4] a_24240_23158# 0.046238f
C1080 ui_in[3] ui_in[2] 5.80246f
C1081 uio_in[4] uio_in[1] 5.22e-19
C1082 uio_in[3] uio_in[2] 8.07582f
C1083 a_12420_37444# VDPWR 0.497771f
C1084 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12310_37398# 3.45e-19
C1085 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.100263f
C1086 tdc_0.diff_gen_0.delay_unit_2_6.in_1 tdc_0.diff_gen_0.delay_unit_2_6.in_2 0.667766f
C1087 input_stage_0.fine_delay_unit_0.in uio_in[5] 0.042742f
C1088 uo_out[2] tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.229249f
C1089 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.499806f
C1090 a_9330_14344# VDPWR 1.1544f
C1091 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 uo_out[3] 3.69e-19
C1092 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.138497f
C1093 a_12310_35116# uo_out[5] 0.098308f
C1094 a_9330_14054# a_9330_15794# 5.08e-20
C1095 a_24240_14314# variable_delay_short_0.variable_delay_unit_1.in 8.82e-20
C1096 ui_in[3] a_25060_11366# 0.002391f
C1097 uo_out[1] tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 1.53e-22
C1098 a_10108_37144# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.007929f
C1099 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_2 0.667766f
C1100 a_24240_21092# a_25060_21092# 0.011184f
C1101 a_15322_7112# a_16292_6702# 0.53267f
C1102 a_12308_26450# VDPWR 1.40782f
C1103 input_stage_0.fine_delay_unit_0.in a_16292_6966# 0.028846f
C1104 input_stage_1.fine_delay_unit_0.in VDPWR 1.5444f
C1105 a_25060_23158# variable_delay_short_0.variable_delay_unit_4.in 8.82e-20
C1106 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_24240_18144# 0.029284f
C1107 ui_in[6] uio_in[3] 9.55e-20
C1108 uio_oe[7] uio_oe[6] 0.170937f
C1109 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 6.93e-19
C1110 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_10108_28016# 0.007929f
C1111 a_12420_28694# a_13254_28694# 0.003413f
C1112 uo_out[1] tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.10528f
C1113 input_stage_1.fine_delay_unit_1.in a_24790_6936# 5.97e-19
C1114 a_16786_5138# VDPWR 0.002853f
C1115 uo_out[6] VDPWR 0.587468f
C1116 tdc_0.start_buffer_0.start_buff tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.001356f
C1117 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_25060_12248# 0.15982f
C1118 a_12310_25988# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 3.84e-19
C1119 variable_delay_dummy_0.variable_delay_unit_1.in a_15680_11634# 0.088132f
C1120 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 8.54e-19
C1121 variable_delay_short_0.out variable_delay_dummy_0.out 1.03552f
C1122 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.747722f
C1123 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 6.79e-20
C1124 tdc_0.diff_gen_0.delay_unit_2_4.in_1 tdc_0.diff_gen_0.delay_unit_2_2.in_1 0.001356f
C1125 a_25060_14314# VDPWR 6.98e-19
C1126 variable_delay_short_0.variable_delay_unit_1.out ui_in[6] 2.67e-19
C1127 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 8.54e-19
C1128 a_24240_12248# VDPWR 1.6584f
C1129 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 a_10108_30298# 0.192064f
C1130 a_25060_12248# variable_delay_short_0.in 7.65e-21
C1131 ui_in[4] a_24240_21092# 6.99e-20
C1132 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.in 0.091118f
C1133 a_12308_28732# a_12310_28270# 0.00595f
C1134 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_12420_28316# 0.013457f
C1135 uio_in[3] variable_delay_dummy_0.out 0.002875f
C1136 uo_out[0] VDPWR 0.587468f
C1137 variable_delay_short_0.variable_delay_unit_5.forward variable_delay_short_0.variable_delay_unit_5.in 0.087283f
C1138 a_12420_35540# VDPWR 0.497547f
C1139 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.283838f
C1140 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 uo_out[5] 0.10528f
C1141 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_13254_23752# 0.010872f
C1142 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_13254_26034# 0.010872f
C1143 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.out 0.002141f
C1144 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 9.61e-20
C1145 input_stage_1.nand_gate_0.out VDPWR 1.47783f
C1146 input_stage_1.fine_delay_unit_1.in input_stage_1.fine_delay_unit_0.in 0.029975f
C1147 a_12420_39726# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.003664f
C1148 ui_in[5] VDPWR 1.43813f
C1149 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_13254_37822# 0.174293f
C1150 a_10108_37144# a_12310_37398# 2.08e-21
C1151 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_13254_23752# 0.005542f
C1152 a_13254_30598# uo_out[3] 0.188081f
C1153 ui_in[5] a_25060_18144# 6.99e-20
C1154 uio_in[0] uio_in[1] 6.17178f
C1155 a_24240_24040# VDPWR 1.65847f
C1156 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_12420_33258# 0.033952f
C1157 a_24240_26106# VDPWR 1.70112f
C1158 a_13254_33258# VDPWR 6.18e-19
C1159 a_12420_33258# uo_out[4] 0.013457f
C1160 tdc_0.start_buffer_0.start_buff a_9330_14054# 1.66e-19
C1161 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[7] 1.09349f
C1162 a_24240_15196# variable_delay_short_0.variable_delay_unit_1.out 0.493816f
C1163 a_15680_15464# VDPWR 1.78268f
C1164 uo_out[7] uo_out[6] 0.856749f
C1165 ui_in[5] variable_delay_short_0.variable_delay_unit_5.out 1.07e-20
C1166 ui_in[3] variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 0.014554f
C1167 a_12308_31014# a_13254_30976# 1.02e-19
C1168 uo_out[1] a_12308_26450# 0.014835f
C1169 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12420_30976# 0.504416f
C1170 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_25060_24040# 0.15982f
C1171 variable_delay_short_0.variable_delay_unit_5.out a_24240_26106# 0.505512f
C1172 variable_delay_short_0.variable_delay_unit_5.out a_24240_24040# 0.071074f
C1173 a_24240_26988# variable_delay_short_0.variable_delay_unit_5.in 7.65e-21
C1174 a_12310_25988# a_13254_26034# 1.02e-19
C1175 ui_in[3] variable_delay_short_0.in 0.052959f
C1176 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 6.79e-20
C1177 a_9330_14344# a_9330_15794# 1.76e-19
C1178 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12308_28732# 0.197073f
C1179 ui_in[3] a_24240_18144# 0.001719f
C1180 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.2373f
C1181 input_stage_0.nand_gate_0.out VDPWR 1.25731f
C1182 uo_out[2] a_13254_28694# 0.005542f
C1183 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_10108_39426# 0.09966f
C1184 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.441213f
C1185 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 uo_out[3] 6.28e-22
C1186 uo_out[5] uo_out[2] 2.26e-21
C1187 uo_out[4] uo_out[3] 1.91867f
C1188 ui_in[1] ui_in[0] 6.25329f
C1189 uio_in[1] uio_in[5] 3.32e-20
C1190 ui_in[4] variable_delay_short_0.variable_delay_unit_4.in 0.507197f
C1191 ui_in[5] a_24240_20210# 0.043085f
C1192 a_13254_37444# VDPWR 6.18e-19
C1193 a_12420_26412# VDPWR 0.497547f
C1194 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.752988f
C1195 ui_in[3] variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 0.014554f
C1196 a_12308_37860# uo_out[6] 0.014835f
C1197 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.192064f
C1198 a_25060_26988# ui_in[3] 0.002391f
C1199 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_10108_37144# 0.09966f
C1200 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.018644f
C1201 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 a_10108_23452# 0.192064f
C1202 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.752988f
C1203 uo_out[0] tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 1.35e-20
C1204 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_10108_32580# 1.06381f
C1205 uo_out[1] uo_out[0] 2.98059f
C1206 a_16292_6966# uio_in[1] 0.022988f
C1207 ui_in[5] uio_in[2] 9.52e-20
C1208 a_24240_14314# variable_delay_short_0.variable_delay_unit_2.in 0.088132f
C1209 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.006183f
C1210 a_12310_25988# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 4.55e-19
C1211 ui_in[5] variable_delay_short_0.variable_delay_unit_3.in 0.506427f
C1212 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en VDPWR 3.87518f
C1213 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en a_15680_12516# 0.029284f
C1214 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 1.24e-19
C1215 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.out 0.12029f
C1216 a_12308_33296# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.36e-21
C1217 a_23820_8460# ui_in[3] 0.010812f
C1218 a_9330_14054# variable_delay_short_0.out 7.21e-19
C1219 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 1.24e-19
C1220 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 a_10108_30298# 0.007929f
C1221 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_12310_28270# 3.45e-19
C1222 uio_in[3] variable_delay_short_0.out 0.036391f
C1223 ui_in[2] variable_delay_short_0.variable_delay_unit_4.in 3.31e-20
C1224 ui_in[0] rst_n 0.031023f
C1225 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en a_24240_23158# 0.11539f
C1226 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.019931f
C1227 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 7.19e-22
C1228 ui_in[5] ui_in[6] 5.05846f
C1229 ui_in[4] ui_in[7] 0.002007f
C1230 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57489f
C1231 input_stage_0.nand_gate_0.out uio_in[2] 6.37e-19
C1232 input_stage_0.fine_delay_unit_0.in uio_in[1] 0.009426f
C1233 variable_delay_dummy_0.variable_delay_unit_1.forward a_16500_14582# 0.054206f
C1234 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en a_25060_26106# 2.39e-19
C1235 a_7140_10670# VDPWR 1.86276f
C1236 a_12420_23752# a_12310_23706# 0.030392f
C1237 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_13254_28316# 0.005542f
C1238 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 8.54e-19
C1239 variable_delay_short_0.variable_delay_unit_1.out variable_delay_short_0.out 0.071795f
C1240 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VDPWR 0.706489f
C1241 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12310_35116# 0.196592f
C1242 a_12420_35162# VDPWR 0.497771f
C1243 uo_out[1] a_12420_26412# 0.013457f
C1244 ui_in[3] variable_delay_short_0.variable_delay_unit_1.in 0.02f
C1245 a_12420_30976# a_13254_30976# 0.003413f
C1246 uio_oe[1] uio_oe[0] 0.170937f
C1247 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en ui_in[3] 0.014554f
C1248 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_12310_37398# 0.014814f
C1249 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 6.08e-20
C1250 variable_delay_short_0.variable_delay_unit_4.out VDPWR 1.3445f
C1251 variable_delay_short_0.variable_delay_unit_5.in VDPWR 2.63444f
C1252 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.747722f
C1253 uio_in[2] variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 2.77e-19
C1254 uio_in[0] a_25060_12248# 0.001909f
C1255 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_12420_32880# 0.003664f
C1256 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12420_28694# 0.033952f
C1257 a_12310_32834# VDPWR 1.42789f
C1258 a_12420_32880# uo_out[4] 0.492009f
C1259 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.99e-19
C1260 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en a_25060_17262# 2.39e-19
C1261 ui_in[7] ui_in[2] 7.13e-19
C1262 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.953579f
C1263 a_24240_11366# a_25060_11366# 0.004142f
C1264 variable_delay_dummy_0.variable_delay_unit_1.out VDPWR 1.61031f
C1265 ui_in[5] variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 1.10207f
C1266 variable_delay_short_0.variable_delay_unit_3.out variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en 0.085059f
C1267 a_16500_11634# variable_delay_dummy_0.in 8.82e-20
C1268 ui_in[4] variable_delay_short_0.variable_delay_unit_5.forward 0.036352f
C1269 variable_delay_dummy_0.variable_delay_unit_1.out a_15680_12516# 0.071074f
C1270 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.871529f
C1271 a_12420_37822# uo_out[6] 0.013457f
C1272 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.283838f
C1273 a_12308_31014# a_12310_30552# 0.00595f
C1274 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_12420_30598# 0.013457f
C1275 a_10108_34862# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.007929f
C1276 a_24790_8050# ui_in[3] 0.00799f
C1277 a_24790_8314# ui_in[1] 4.3e-19
C1278 a_12310_32834# tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 1.15e-21
C1279 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_4.out 0.071795f
C1280 variable_delay_short_0.variable_delay_unit_5.out variable_delay_short_0.variable_delay_unit_5.in 0.499092f
C1281 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 a_10108_23452# 0.007929f
C1282 ui_in[1] VDPWR 0.00509f
C1283 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.283838f
C1284 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.871529f
C1285 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.953579f
C1286 uo_out[0] tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 3.69e-19
C1287 uo_out[2] a_12310_28270# 0.098308f
C1288 ui_in[3] variable_delay_short_0.variable_delay_unit_2.out 0.040959f
C1289 a_15322_7112# input_stage_0.nand_gate_0.out 3.78e-19
C1290 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VDPWR 0.706518f
C1291 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.231672f
C1292 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_2.in 0.09141f
C1293 a_12308_35578# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.36e-21
C1294 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 4.28924f
C1295 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.499806f
C1296 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 VDPWR 5.07283f
C1297 a_9330_14344# variable_delay_short_0.out 3.54e-19
C1298 tdc_0.diff_gen_0.delay_unit_2_1.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.667766f
C1299 a_12420_26034# VDPWR 0.497771f
C1300 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 8.54e-19
C1301 variable_delay_short_0.variable_delay_unit_5.out ui_in[1] 0.001119f
C1302 a_9330_14344# a_9330_14054# 0.083149f
C1303 variable_delay_dummy_0.variable_delay_unit_1.out a_15680_14582# 0.505512f
C1304 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.231672f
C1305 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 8.54e-19
C1306 a_12308_33296# a_12420_33258# 0.030083f
C1307 a_12308_31014# VDPWR 1.40782f
C1308 ui_in[4] a_24240_26988# 0.005915f
C1309 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_10108_28016# 1.06381f
C1310 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 0.752988f
C1311 uio_in[0] ui_in[3] 0.014973f
C1312 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 0.132512f
C1313 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.003768f
C1314 variable_delay_short_0.variable_delay_unit_5.forward ui_in[2] 1.68e-20
C1315 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.441213f
C1316 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 uo_out[4] 3.69e-19
C1317 tdc_0.diff_gen_0.delay_unit_2_1.in_1 VDPWR 4.44048f
C1318 a_12310_37398# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 3.84e-19
C1319 a_25060_23158# VDPWR 6.98e-19
C1320 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en variable_delay_dummy_0.out 0.12022f
C1321 ui_in[3] a_25060_20210# 0.002391f
C1322 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12308_31014# 0.197073f
C1323 input_stage_1.fine_delay_unit_1.in ui_in[1] 0.039118f
C1324 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en VDPWR 2.77611f
C1325 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_12310_28270# 3.84e-19
C1326 uio_in[5] ua[0] 0.081349f
C1327 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 1.24e-19
C1328 a_12420_28316# a_12310_28270# 0.030392f
C1329 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 uo_out[3] 0.20241f
C1330 a_13254_24130# VDPWR 6.18e-19
C1331 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 0.192064f
C1332 variable_delay_short_0.out a_24240_12248# 0.493816f
C1333 uo_out[2] tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.10528f
C1334 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_4.in 0.09141f
C1335 a_12308_26450# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.197073f
C1336 ui_in[2] ui_in[0] 0.001501f
C1337 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en a_24240_11366# 0.11539f
C1338 variable_delay_dummy_0.variable_delay_unit_1.in variable_delay_dummy_0.in 0.08442f
C1339 ui_in[3] a_25060_17262# 0.002391f
C1340 ui_in[3] variable_delay_short_0.variable_delay_unit_3.out 0.040959f
C1341 a_16500_11634# VDPWR 0.160518f
C1342 a_12310_23706# a_13254_23752# 1.02e-19
C1343 a_24240_11366# variable_delay_short_0.in 8.82e-20
C1344 ui_in[6] variable_delay_short_0.variable_delay_unit_5.in 0.001598f
C1345 variable_delay_dummy_0.out a_7140_10670# 0.087271f
C1346 tdc_0.start_buffer_0.start_delay a_9330_13764# 1.56e-19
C1347 a_12310_35116# tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.15e-21
C1348 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 VDPWR 5.07283f
C1349 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 6.93e-19
C1350 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VDPWR 2.55561f
C1351 ui_in[7] variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en 9.38e-20
C1352 variable_delay_short_0.variable_delay_unit_1.out a_25060_14314# 0.222585f
C1353 a_13254_35162# VDPWR 6.18e-19
C1354 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_10108_23452# 0.09966f
C1355 variable_delay_short_0.variable_delay_unit_1.out a_24240_12248# 0.071074f
C1356 a_12308_35578# uo_out[6] 6.49e-20
C1357 uo_out[0] tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.10528f
C1358 a_23820_7082# a_24790_6672# 0.53267f
C1359 uo_out[1] a_12420_26034# 0.492009f
C1360 input_stage_1.fine_delay_unit_0.in a_24790_6936# 0.028846f
C1361 ui_in[3] variable_delay_short_0.variable_delay_unit_2.in 0.02f
C1362 uo_out[0] uio_in[7] 0.073214f
C1363 a_16292_6702# input_stage_0.nand_gate_0.out 5.26e-20
C1364 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.019931f
C1365 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 VDPWR 2.57093f
C1366 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.138497f
C1367 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 6.93e-19
C1368 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.138497f
C1369 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.019931f
C1370 a_25060_21092# VDPWR 0.001468f
C1371 uo_out[0] tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 6.28e-22
C1372 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_12420_28316# 0.003664f
C1373 a_12420_40104# a_13254_40104# 0.003413f
C1374 a_13254_32880# uo_out[4] 0.188081f
C1375 a_13254_28694# VDPWR 6.18e-19
C1376 input_stage_0.fine_delay_unit_0.in ua[0] 4.88e-20
C1377 tdc_0.start_buffer_0.start_buff a_7140_10670# 0.684455f
C1378 a_12308_35578# a_12420_35540# 0.030083f
C1379 uo_out[5] VDPWR 0.587468f
C1380 variable_delay_dummy_0.variable_delay_unit_1.out variable_delay_dummy_0.out 0.071795f
C1381 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.2373f
C1382 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en a_15680_15464# 0.029284f
C1383 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.196592f
C1384 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_3.in 7.91e-21
C1385 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_13254_30598# 0.005542f
C1386 a_12420_37444# uo_out[6] 0.492009f
C1387 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 1.24e-19
C1388 variable_delay_short_0.variable_delay_unit_4.out variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 0.085059f
C1389 variable_delay_short_0.variable_delay_unit_5.in variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en 7.91e-21
C1390 uio_oe[6] uio_oe[5] 0.170937f
C1391 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_13254_37822# 0.012202f
C1392 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 1.24e-19
C1393 a_12420_30976# VDPWR 0.497547f
C1394 a_12310_39680# tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.45e-19
C1395 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.871529f
C1396 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 0.283838f
C1397 ui_in[4] VDPWR 1.64573f
C1398 uo_out[7] tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.203149f
C1399 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.99e-19
C1400 a_25060_15196# ui_in[3] 0.002391f
C1401 uio_in[7] uio_in[6] 0.073214f
C1402 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 uo_out[4] 6.28e-22
C1403 uio_in[5] a_15680_11634# 0.002316f
C1404 uio_in[2] a_16500_11634# 3.05e-20
C1405 a_12310_37398# tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 4.55e-19
C1406 a_24790_6936# input_stage_1.nand_gate_0.out 4.47e-20
C1407 a_13254_26034# VDPWR 6.18e-19
C1408 variable_delay_short_0.out variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 2.24e-20
C1409 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_12420_30976# 0.033952f
C1410 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en ui_in[6] 9.38e-20
C1411 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_12310_28270# 4.55e-19
C1412 a_10108_32580# a_12310_32834# 2.08e-21
C1413 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_13254_33258# 0.174293f
C1414 variable_delay_dummy_0.variable_delay_unit_1.in VDPWR 3.21199f
C1415 ui_in[4] variable_delay_short_0.variable_delay_unit_5.out 0.047464f
C1416 uio_in[3] variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.00127f
C1417 a_10108_25734# tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.007929f
C1418 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.752988f
C1419 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.132512f
C1420 variable_delay_dummy_0.variable_delay_unit_1.in a_15680_12516# 0.020173f
C1421 uo_out[1] tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 1.35e-20
C1422 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_12308_40142# 0.162625f
C1423 variable_delay_short_0.variable_delay_unit_5.forward variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en 7.91e-21
C1424 ui_in[7] uio_in[4] 3.77e-20
C1425 a_12420_26412# tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.033952f
C1426 uo_out[7] uo_out[5] 1.56e-19
C1427 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12310_37398# 6.08e-20
C1428 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12308_40142# 2.36e-21
C1429 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en 0.002365f
C1430 a_9330_15504# tdc_0.diff_gen_0.delay_unit_2_1.in_1 8.59e-20
C1431 variable_delay_short_0.variable_delay_unit_1.in a_24240_11366# 0.088132f
C1432 a_12308_37860# tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 7.19e-22
C1433 a_25060_21092# variable_delay_short_0.variable_delay_unit_3.in 7.65e-21
C1434 a_24240_21092# variable_delay_short_0.variable_delay_unit_3.out 0.493816f
C1435 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_12308_37860# 0.162625f
C1436 a_24790_8314# ui_in[2] 0.024917f
C1437 ui_in[2] VDPWR 0.001157f
C1438 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_12308_28732# 7.19e-22
C1439 a_12308_31014# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.36e-21
C1440 a_12310_28270# a_13254_28316# 1.02e-19
C1441 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 a_12310_30552# 3.84e-19
C1442 a_9330_15214# a_9330_14924# 0.083149f
C1443 input_stage_1.fine_delay_unit_0.in input_stage_1.nand_gate_0.out 0.062526f
C1444 ui_in[2] a_25060_18144# 3.98e-20
C1445 a_12310_23706# VDPWR 1.42748f
C1446 tdc_0.diff_gen_0.delay_unit_2_2.in_2 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.311186f
C1447 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 VDPWR 3.23832f
C1448 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.018644f
C1449 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 a_10108_32580# 0.192064f
C1450 uo_out[4] uo_out[2] 1.56e-19
C1451 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en a_24240_15196# 0.029284f
C1452 ui_in[7] variable_delay_short_0.variable_delay_unit_1.in 0.506369f
C1453 a_15680_14582# variable_delay_dummy_0.variable_delay_unit_1.in 8.82e-20
C1454 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.441213f
C1455 a_12420_37444# a_13254_37444# 0.003413f
C1456 variable_delay_short_0.variable_delay_unit_5.out ui_in[2] 0.002549f
C1457 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_10108_30298# 1.06381f
C1458 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.871529f
C1459 a_12420_40104# VDPWR 0.497547f
C1460 a_25060_11366# VDPWR 6.98e-19
C1461 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 4.28924f
C1462 tdc_0.start_buffer_0.start_buff tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.751615f
C1463 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.018644f
C1464 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.441213f
C1465 variable_delay_dummy_0.out a_16500_11634# 0.222585f
C1466 a_24240_26988# a_25060_26988# 0.011184f
C1467 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 1.17e-19
C1468 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 a_12308_33296# 5.04e-20
C1469 tdc_0.vernier_delay_line_0.start_pos tdc_0.vernier_delay_line_0.start_neg 0.688629f
C1470 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 VDPWR 5.07283f
C1471 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.231672f
C1472 variable_delay_short_0.variable_delay_unit_4.in a_25060_20210# 0.054206f
C1473 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.747722f
C1474 uio_in[2] variable_delay_dummy_0.variable_delay_unit_1.in 1.1e-20
C1475 uo_out[1] a_13254_26034# 0.188081f
C1476 a_12420_30598# a_12310_30552# 0.030392f
C1477 tdc_0.vernier_delay_line_0.start_neg tdc_0.diff_gen_0.delay_unit_2_6.in_2 0.036472f
C1478 input_stage_1.fine_delay_unit_1.in ui_in[2] 0.010002f
C1479 ui_in[7] variable_delay_short_0.variable_delay_unit_2.out 0.043504f
C1480 a_12308_26450# a_12420_26412# 0.030083f
C1481 variable_delay_dummy_0.variable_delay_unit_1.out uio_in[3] 3.5e-20
C1482 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.138497f
C1483 input_stage_0.nand_gate_0.out a_16786_5138# 0.355469f
C1484 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.019931f
C1485 ui_in[1] variable_delay_short_0.out 0.001119f
C1486 uio_in[0] a_24240_11366# 0.042718f
C1487 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 4.53e-19
C1488 tdc_0.diff_gen_0.delay_unit_2_2.in_1 tdc_0.diff_gen_0.delay_unit_2_1.in_1 0.756572f
C1489 a_12310_28270# VDPWR 1.42789f
C1490 ui_in[4] ui_in[6] 0.002613f
C1491 variable_delay_short_0.variable_delay_unit_4.in variable_delay_short_0.variable_delay_unit_3.out 0.235667f
C1492 a_24240_14314# ui_in[3] 0.001719f
C1493 a_10108_34862# a_12310_35116# 2.08e-21
C1494 variable_delay_dummy_0.in a_16292_8344# 7.3e-20
C1495 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13254_35540# 0.174293f
C1496 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en variable_delay_dummy_0.variable_delay_unit_1.out 0.12029f
C1497 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en variable_delay_short_0.variable_delay_unit_5.forward 0.794183f
C1498 ui_in[5] a_24240_24040# 2.89e-20
C1499 a_13254_37444# uo_out[6] 0.188081f
C1500 ui_in[2] variable_delay_short_0.variable_delay_unit_3.in 3.31e-20
C1501 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en a_25060_21092# 0.15982f
C1502 a_12310_35116# tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 3.84e-19
C1503 a_12420_40104# uo_out[7] 0.013457f
C1504 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12310_37398# 0.164402f
C1505 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 a_12310_23706# 3.84e-19
C1506 a_9330_14924# a_9330_14634# 0.083149f
C1507 ui_in[7] uio_in[0] 9.98875f
C1508 a_12310_30552# tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.15e-21
C1509 a_12420_30598# VDPWR 0.497771f
C1510 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.283838f
C1511 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.871529f
C1512 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_12310_32834# 0.196592f
C1513 a_12310_35116# a_12308_33296# 0.005984f
C1514 uo_out[1] tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 3.69e-19
C1515 ua[1] VGND 0.146962f
C1516 ua[2] VGND 0.146962f
C1517 ua[3] VGND 0.146962f
C1518 ua[4] VGND 0.146962f
C1519 ua[5] VGND 0.146962f
C1520 ua[6] VGND 0.146962f
C1521 ua[7] VGND 0.146962f
C1522 ena VGND 0.070385f
C1523 clk VGND 0.042875f
C1524 rst_n VGND 0.042875f
C1525 uio_in[6] VGND 0.071255f
C1526 uio_in[7] VGND 0.071255f
C1527 uio_out[0] VGND 0.136988f
C1528 uio_out[1] VGND 0.136988f
C1529 uio_out[2] VGND 0.137343f
C1530 uio_out[3] VGND 0.137343f
C1531 uio_out[4] VGND 0.137343f
C1532 uio_out[5] VGND 0.137343f
C1533 uio_out[6] VGND 0.137343f
C1534 uio_out[7] VGND 0.137343f
C1535 uio_oe[0] VGND 0.137343f
C1536 uio_oe[1] VGND 0.137343f
C1537 uio_oe[2] VGND 0.137343f
C1538 uio_oe[3] VGND 0.137339f
C1539 uio_oe[4] VGND 0.137343f
C1540 uio_oe[5] VGND 0.137343f
C1541 uio_oe[6] VGND 0.137343f
C1542 uio_oe[7] VGND 0.289256f
C1543 ua[0] VGND 11.616f
C1544 uio_in[5] VGND 15.11678f
C1545 ui_in[0] VGND 14.124138f
C1546 ui_in[1] VGND 12.519405f
C1547 uio_in[1] VGND 15.046968f
C1548 uio_in[2] VGND 15.199068f
C1549 ui_in[2] VGND 11.54435f
C1550 ui_in[3] VGND 12.04699f
C1551 uio_in[3] VGND 14.21004f
C1552 uio_in[4] VGND 14.381983f
C1553 uio_in[0] VGND 15.490564f
C1554 ui_in[7] VGND 15.539585f
C1555 ui_in[6] VGND 12.882964f
C1556 ui_in[5] VGND 10.864614f
C1557 ui_in[4] VGND 9.591749f
C1558 uo_out[0] VGND 8.491008f
C1559 uo_out[1] VGND 8.284716f
C1560 uo_out[2] VGND 7.409694f
C1561 uo_out[3] VGND 5.486512f
C1562 uo_out[4] VGND 3.7559f
C1563 uo_out[5] VGND 3.29391f
C1564 uo_out[6] VGND 2.83951f
C1565 uo_out[7] VGND 2.66217f
C1566 VDPWR VGND 0.359394p
C1567 a_25284_5108# VGND 0.372398f
C1568 a_16786_5138# VGND 0.37196f
C1569 input_stage_1.nand_gate_0.out VGND 0.885485f
C1570 input_stage_0.nand_gate_0.out VGND 0.872828f
C1571 a_24790_6672# VGND 0.387205f
C1572 a_24790_6936# VGND 0.612975f
C1573 input_stage_1.fine_delay_unit_0.in VGND 1.83045f
C1574 a_23820_7082# VGND 0.731446f
C1575 a_16292_6702# VGND 0.387205f
C1576 a_16292_6966# VGND 0.612975f
C1577 input_stage_0.fine_delay_unit_0.in VGND 1.8013f
C1578 a_15322_7112# VGND 0.731446f
C1579 a_24790_8050# VGND 0.387205f
C1580 a_24790_8314# VGND 0.612975f
C1581 input_stage_1.fine_delay_unit_1.in VGND 1.68519f
C1582 a_23820_8460# VGND 0.739963f
C1583 a_16292_8080# VGND 0.387205f
C1584 a_16292_8344# VGND 0.612975f
C1585 input_stage_0.fine_delay_unit_1.in VGND 1.67858f
C1586 a_15322_8490# VGND 0.739963f
C1587 variable_delay_short_0.in VGND 1.97381f
C1588 variable_delay_dummy_0.in VGND 1.96449f
C1589 a_25060_11366# VGND 0.71648f
C1590 a_24240_11366# VGND 0.037888f
C1591 a_16500_11634# VGND 0.71648f
C1592 a_15680_11634# VGND 0.037888f
C1593 a_7140_10670# VGND 1.49885f
C1594 a_25060_12248# VGND 0.717347f
C1595 a_24240_12248# VGND 0.043128f
C1596 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en VGND 2.516856f
C1597 variable_delay_dummy_0.out VGND 5.71113f
C1598 a_16500_12516# VGND 0.717347f
C1599 a_15680_12516# VGND 0.043128f
C1600 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en VGND 2.851508f
C1601 variable_delay_short_0.variable_delay_unit_1.in VGND 3.604031f
C1602 variable_delay_short_0.out VGND 8.859031f
C1603 variable_delay_dummy_0.variable_delay_unit_1.in VGND 4.168124f
C1604 a_9330_13764# VGND 0.629875f
C1605 a_25060_14314# VGND 0.71648f
C1606 a_24240_14314# VGND 0.037888f
C1607 a_9330_14054# VGND 0.622523f
C1608 tdc_0.start_buffer_0.start_delay VGND 3.694501f
C1609 tdc_0.start_buffer_0.start_buff VGND 5.257338f
C1610 a_16500_14582# VGND 0.71648f
C1611 a_15680_14582# VGND 0.037888f
C1612 variable_delay_dummy_0.variable_delay_unit_1.forward VGND 2.636476f
C1613 a_9330_14344# VGND 0.622523f
C1614 a_9330_14634# VGND 0.622248f
C1615 variable_delay_short_0.variable_delay_unit_1.out VGND 2.21957f
C1616 a_25060_15196# VGND 0.717347f
C1617 a_24240_15196# VGND 0.043128f
C1618 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en VGND 2.517556f
C1619 a_9330_14924# VGND 0.622523f
C1620 variable_delay_dummy_0.variable_delay_unit_1.out VGND 2.29732f
C1621 a_16500_15464# VGND 0.784074f
C1622 a_15680_15464# VGND 0.114203f
C1623 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en VGND 2.963248f
C1624 a_9330_15214# VGND 0.622289f
C1625 a_9330_15504# VGND 0.622536f
C1626 tdc_0.diff_gen_0.delay_unit_2_1.in_2 VGND 3.077349f
C1627 tdc_0.diff_gen_0.delay_unit_2_1.in_1 VGND 2.012721f
C1628 variable_delay_short_0.variable_delay_unit_2.in VGND 3.604041f
C1629 a_9330_15794# VGND 1.49187f
C1630 tdc_0.diff_gen_0.delay_unit_2_2.in_2 VGND 3.163373f
C1631 tdc_0.diff_gen_0.delay_unit_2_2.in_1 VGND 2.006561f
C1632 a_25060_17262# VGND 0.71648f
C1633 a_24240_17262# VGND 0.037888f
C1634 variable_delay_short_0.variable_delay_unit_2.out VGND 2.21957f
C1635 a_25060_18144# VGND 0.717347f
C1636 a_24240_18144# VGND 0.043128f
C1637 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en VGND 2.517556f
C1638 tdc_0.diff_gen_0.delay_unit_2_3.in_2 VGND 3.077369f
C1639 tdc_0.diff_gen_0.delay_unit_2_3.in_1 VGND 2.006501f
C1640 variable_delay_short_0.variable_delay_unit_3.in VGND 3.604041f
C1641 tdc_0.diff_gen_0.delay_unit_2_4.in_2 VGND 3.163433f
C1642 tdc_0.diff_gen_0.delay_unit_2_4.in_1 VGND 2.006681f
C1643 a_25060_20210# VGND 0.71648f
C1644 a_24240_20210# VGND 0.037888f
C1645 tdc_0.diff_gen_0.delay_unit_2_5.in_2 VGND 3.163143f
C1646 variable_delay_short_0.variable_delay_unit_3.out VGND 2.21957f
C1647 a_25060_21092# VGND 0.717347f
C1648 a_24240_21092# VGND 0.043128f
C1649 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en VGND 2.517556f
C1650 tdc_0.diff_gen_0.delay_unit_2_6.in_2 VGND 3.083859f
C1651 tdc_0.diff_gen_0.delay_unit_2_6.in_1 VGND 2.070971f
C1652 variable_delay_short_0.variable_delay_unit_4.in VGND 3.604041f
C1653 a_25060_23158# VGND 0.71648f
C1654 a_24240_23158# VGND 0.037888f
C1655 variable_delay_short_0.variable_delay_unit_4.out VGND 2.21957f
C1656 a_25060_24040# VGND 0.717347f
C1657 a_24240_24040# VGND 0.043128f
C1658 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en VGND 2.517556f
C1659 a_13254_23752# VGND 0.190873f
C1660 a_12310_23706# VGND 0.838649f
C1661 a_12420_23752# VGND 0.024712f
C1662 a_13254_24130# VGND 0.192269f
C1663 a_12420_24130# VGND 0.023462f
C1664 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VGND 0.583709f
C1665 a_12308_24168# VGND 0.823328f
C1666 a_10108_23452# VGND 0.354057f
C1667 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 VGND 6.034074f
C1668 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 VGND 7.095738f
C1669 tdc_0.vernier_delay_line_0.start_neg VGND 3.594784f
C1670 tdc_0.vernier_delay_line_0.start_pos VGND 2.750328f
C1671 variable_delay_short_0.variable_delay_unit_5.in VGND 3.860429f
C1672 a_25060_26106# VGND 0.71648f
C1673 a_24240_26106# VGND 0.037888f
C1674 variable_delay_short_0.variable_delay_unit_5.forward VGND 2.636476f
C1675 a_13254_26034# VGND 0.190624f
C1676 a_12310_25988# VGND 0.829382f
C1677 a_12420_26034# VGND 0.024712f
C1678 a_13254_26412# VGND 0.192129f
C1679 a_12420_26412# VGND 0.023462f
C1680 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VGND 0.583105f
C1681 a_12308_26450# VGND 0.823144f
C1682 variable_delay_short_0.variable_delay_unit_5.out VGND 2.29732f
C1683 a_25060_26988# VGND 0.784074f
C1684 a_24240_26988# VGND 0.114203f
C1685 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en VGND 2.963248f
C1686 a_10108_25734# VGND 0.354057f
C1687 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1688 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1689 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 VGND 6.192364f
C1690 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 VGND 5.851951f
C1691 a_13254_28316# VGND 0.190624f
C1692 a_12310_28270# VGND 0.829382f
C1693 a_12420_28316# VGND 0.024712f
C1694 a_13254_28694# VGND 0.192129f
C1695 a_12420_28694# VGND 0.023462f
C1696 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VGND 0.583105f
C1697 a_12308_28732# VGND 0.823144f
C1698 a_10108_28016# VGND 0.354057f
C1699 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1700 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1701 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 VGND 6.192265f
C1702 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 VGND 5.68077f
C1703 a_13254_30598# VGND 0.190624f
C1704 a_12310_30552# VGND 0.829382f
C1705 a_12420_30598# VGND 0.024712f
C1706 a_13254_30976# VGND 0.192129f
C1707 a_12420_30976# VGND 0.023462f
C1708 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VGND 0.583105f
C1709 a_12308_31014# VGND 0.823144f
C1710 a_10108_30298# VGND 0.354057f
C1711 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1712 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1713 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 VGND 6.192265f
C1714 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 VGND 5.68077f
C1715 a_13254_32880# VGND 0.190624f
C1716 a_12310_32834# VGND 0.829382f
C1717 a_12420_32880# VGND 0.024712f
C1718 a_13254_33258# VGND 0.192129f
C1719 a_12420_33258# VGND 0.023462f
C1720 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VGND 0.583105f
C1721 a_12308_33296# VGND 0.823144f
C1722 a_10108_32580# VGND 0.354057f
C1723 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1724 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1725 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 VGND 6.021708f
C1726 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 VGND 5.489025f
C1727 a_13254_35162# VGND 0.190624f
C1728 a_12310_35116# VGND 0.829382f
C1729 a_12420_35162# VGND 0.024712f
C1730 a_13254_35540# VGND 0.192129f
C1731 a_12420_35540# VGND 0.023462f
C1732 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VGND 0.583105f
C1733 a_12308_35578# VGND 0.823144f
C1734 a_10108_34862# VGND 0.354057f
C1735 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1736 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1737 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 VGND 6.021708f
C1738 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 VGND 5.489025f
C1739 a_13254_37444# VGND 0.190624f
C1740 a_12310_37398# VGND 0.829382f
C1741 a_12420_37444# VGND 0.024712f
C1742 a_13254_37822# VGND 0.192129f
C1743 a_12420_37822# VGND 0.023462f
C1744 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VGND 0.583105f
C1745 a_12308_37860# VGND 0.823144f
C1746 a_10108_37144# VGND 0.354057f
C1747 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 VGND 6.032664f
C1748 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 VGND 6.447248f
C1749 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 VGND 6.192265f
C1750 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 VGND 5.68077f
C1751 a_13254_39726# VGND 0.190624f
C1752 a_12310_39680# VGND 0.829382f
C1753 a_12420_39726# VGND 0.024712f
C1754 a_13254_40104# VGND 0.192129f
C1755 a_12420_40104# VGND 0.023462f
C1756 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VGND 0.583308f
C1757 a_12308_40142# VGND 0.830326f
C1758 a_10108_39426# VGND 0.354057f
C1759 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VGND 6.505114f
C1760 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 VGND 6.446748f
C1761 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 VGND 6.192265f
C1762 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 VGND 5.68077f
C1763 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1 VGND 0.974288f
C1764 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_2 VGND 1.24637f
C1765 uio_in[2].t0 VGND 0.083134f
C1766 uio_in[2].n0 VGND 7.1868f
C1767 ui_in[1].t0 VGND 0.062351f
C1768 ui_in[1].n0 VGND 4.87703f
C1769 uio_in[5].t0 VGND 0.026624f
C1770 uio_in[5].t1 VGND 0.035892f
C1771 uio_in[5].n0 VGND 0.039941f
C1772 uio_in[5].n1 VGND 2.89986f
C1773 uio_in[4].t0 VGND 0.084602f
C1774 uio_in[4].n0 VGND 6.89354f
C1775 uio_in[1].t0 VGND 0.064466f
C1776 uio_in[1].n0 VGND 6.45166f
C1777 ui_in[3].t0 VGND 0.046163f
C1778 ui_in[3].n0 VGND 3.40417f
C1779 variable_delay_short_0.variable_delay_unit_1.in.t4 VGND 0.017058f
C1780 variable_delay_short_0.variable_delay_unit_1.in.t5 VGND 0.044984f
C1781 variable_delay_short_0.variable_delay_unit_1.in.n0 VGND 0.04731f
C1782 variable_delay_short_0.variable_delay_unit_1.in.t0 VGND 0.033139f
C1783 variable_delay_short_0.variable_delay_unit_1.in.t1 VGND 0.105354f
C1784 variable_delay_short_0.variable_delay_unit_1.in.n1 VGND 0.255341f
C1785 variable_delay_short_0.variable_delay_unit_1.in.t2 VGND 0.042943f
C1786 variable_delay_short_0.variable_delay_unit_1.in.t3 VGND 0.013862f
C1787 variable_delay_short_0.variable_delay_unit_1.in.n2 VGND 0.045161f
C1788 variable_delay_short_0.variable_delay_unit_1.in.n3 VGND 0.418008f
C1789 variable_delay_short_0.variable_delay_unit_2.in.t4 VGND 0.017058f
C1790 variable_delay_short_0.variable_delay_unit_2.in.t5 VGND 0.044984f
C1791 variable_delay_short_0.variable_delay_unit_2.in.n0 VGND 0.04731f
C1792 variable_delay_short_0.variable_delay_unit_2.in.t1 VGND 0.033139f
C1793 variable_delay_short_0.variable_delay_unit_2.in.t0 VGND 0.105354f
C1794 variable_delay_short_0.variable_delay_unit_2.in.n1 VGND 0.255341f
C1795 variable_delay_short_0.variable_delay_unit_2.in.t2 VGND 0.042943f
C1796 variable_delay_short_0.variable_delay_unit_2.in.t3 VGND 0.013862f
C1797 variable_delay_short_0.variable_delay_unit_2.in.n2 VGND 0.045161f
C1798 variable_delay_short_0.variable_delay_unit_2.in.n3 VGND 0.418008f
C1799 a_10108_37672.t3 VGND 0.059028f
C1800 a_10108_37672.t2 VGND 0.059028f
C1801 a_10108_37672.t5 VGND 0.059028f
C1802 a_10108_37672.n0 VGND 0.136068f
C1803 a_10108_37672.t0 VGND 0.059028f
C1804 a_10108_37672.t1 VGND 0.059028f
C1805 a_10108_37672.n1 VGND 0.139449f
C1806 a_10108_37672.n2 VGND 1.11221f
C1807 a_10108_37672.n3 VGND 0.258102f
C1808 a_10108_37672.t4 VGND 0.059028f
C1809 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 VGND 0.930597f
C1810 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.765644f
C1811 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.087567f
C1812 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C1813 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C1814 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C1815 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.054262f
C1816 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C1817 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.115417f
C1818 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.089004f
C1819 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C1820 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C1821 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.041221f
C1822 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.095888f
C1823 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C1824 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.108461f
C1825 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.202442f
C1826 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 VGND 0.748416f
C1827 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C1828 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.041341f
C1829 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.096169f
C1830 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C1831 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.089265f
C1832 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.083414f
C1833 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C1834 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.202074f
C1835 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.087824f
C1836 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C1837 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C1838 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.200787f
C1839 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C1840 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.054421f
C1841 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C1842 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C1843 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.107523f
C1844 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C1845 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C1846 ui_in[0].t0 VGND 0.028496f
C1847 ui_in[0].n0 VGND 2.53887f
C1848 uio_in[3].t0 VGND 0.07563f
C1849 uio_in[3].n0 VGND 7.04584f
C1850 uo_out[2].t5 VGND 0.01472f
C1851 uo_out[2].t4 VGND 0.04976f
C1852 uo_out[2].n0 VGND 0.040339f
C1853 uo_out[2].t2 VGND 0.028671f
C1854 uo_out[2].t1 VGND 0.028671f
C1855 uo_out[2].n1 VGND 0.060931f
C1856 uo_out[2].n2 VGND 0.265829f
C1857 uo_out[2].t0 VGND 0.009557f
C1858 uo_out[2].t3 VGND 0.009557f
C1859 uo_out[2].n3 VGND 0.020748f
C1860 uo_out[2].n4 VGND 0.070592f
C1861 uo_out[2].n5 VGND 1.57081f
C1862 uo_out[1].t5 VGND 0.015076f
C1863 uo_out[1].t4 VGND 0.050965f
C1864 uo_out[1].n0 VGND 0.041315f
C1865 uo_out[1].t0 VGND 0.029365f
C1866 uo_out[1].t3 VGND 0.029365f
C1867 uo_out[1].n1 VGND 0.062406f
C1868 uo_out[1].n2 VGND 0.272264f
C1869 uo_out[1].t2 VGND 0.009788f
C1870 uo_out[1].t1 VGND 0.009788f
C1871 uo_out[1].n3 VGND 0.02125f
C1872 uo_out[1].n4 VGND 0.072301f
C1873 uo_out[1].n5 VGND 1.84327f
C1874 ui_in[2].t0 VGND 0.055937f
C1875 ui_in[2].n0 VGND 4.70026f
C1876 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t2 VGND 0.020532f
C1877 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t0 VGND 0.020532f
C1878 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n0 VGND 0.048092f
C1879 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t4 VGND 0.061597f
C1880 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t5 VGND 0.061597f
C1881 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n1 VGND 0.125485f
C1882 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n2 VGND 0.522094f
C1883 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t1 VGND 0.075157f
C1884 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.t3 VGND 0.227425f
C1885 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n3 VGND 0.55466f
C1886 tdc_0.vernier_delay_line_0.delay_unit_2_0.out_1.n4 VGND 0.283681f
C1887 variable_delay_dummy_0.variable_delay_unit_1.forward.t3 VGND 0.025654f
C1888 variable_delay_dummy_0.variable_delay_unit_1.forward.t2 VGND 0.067654f
C1889 variable_delay_dummy_0.variable_delay_unit_1.forward.n0 VGND 0.071153f
C1890 variable_delay_dummy_0.variable_delay_unit_1.forward.t0 VGND 0.04984f
C1891 variable_delay_dummy_0.variable_delay_unit_1.forward.t1 VGND 0.15845f
C1892 variable_delay_dummy_0.variable_delay_unit_1.forward.n1 VGND 0.384027f
C1893 variable_delay_dummy_0.variable_delay_unit_1.forward.n2 VGND 0.628675f
C1894 variable_delay_dummy_0.variable_delay_unit_1.in.t5 VGND 0.025993f
C1895 variable_delay_dummy_0.variable_delay_unit_1.in.t4 VGND 0.068546f
C1896 variable_delay_dummy_0.variable_delay_unit_1.in.n0 VGND 0.072091f
C1897 variable_delay_dummy_0.variable_delay_unit_1.in.t0 VGND 0.050497f
C1898 variable_delay_dummy_0.variable_delay_unit_1.in.t1 VGND 0.160539f
C1899 variable_delay_dummy_0.variable_delay_unit_1.in.n1 VGND 0.389091f
C1900 variable_delay_dummy_0.variable_delay_unit_1.in.t3 VGND 0.065437f
C1901 variable_delay_dummy_0.variable_delay_unit_1.in.t2 VGND 0.021123f
C1902 variable_delay_dummy_0.variable_delay_unit_1.in.n2 VGND 0.068816f
C1903 variable_delay_dummy_0.variable_delay_unit_1.in.n3 VGND 0.636965f
C1904 a_10108_33108.t1 VGND 0.059028f
C1905 a_10108_33108.t0 VGND 0.059028f
C1906 a_10108_33108.t2 VGND 0.059028f
C1907 a_10108_33108.n0 VGND 0.136068f
C1908 a_10108_33108.t5 VGND 0.059028f
C1909 a_10108_33108.t4 VGND 0.059028f
C1910 a_10108_33108.n1 VGND 0.139449f
C1911 a_10108_33108.n2 VGND 1.11221f
C1912 a_10108_33108.n3 VGND 0.258102f
C1913 a_10108_33108.t3 VGND 0.059028f
C1914 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 VGND 0.09757f
C1915 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 VGND 0.030153f
C1916 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 VGND 0.265657f
C1917 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 VGND 0.039259f
C1918 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 VGND 0.012524f
C1919 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 VGND 0.027534f
C1920 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 VGND 0.039259f
C1921 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 VGND 0.012524f
C1922 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 VGND 0.027357f
C1923 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 VGND 0.008823f
C1924 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 VGND 0.039259f
C1925 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 VGND 0.012524f
C1926 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 VGND 0.027534f
C1927 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 VGND 0.039259f
C1928 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 VGND 0.012524f
C1929 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 VGND 0.027357f
C1930 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 VGND 0.008728f
C1931 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 VGND 0.135162f
C1932 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 VGND 0.046129f
C1933 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 VGND 0.046129f
C1934 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 VGND 0.054044f
C1935 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 VGND 0.046129f
C1936 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 VGND 0.046129f
C1937 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 VGND 0.0538f
C1938 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 VGND 0.495704f
C1939 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 VGND 0.119944f
C1940 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 VGND 0.025758f
C1941 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 VGND 0.025758f
C1942 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 VGND 0.055083f
C1943 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 VGND 0.008586f
C1944 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 VGND 0.008586f
C1945 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 VGND 0.01864f
C1946 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 VGND 0.221512f
C1947 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 VGND 0.09757f
C1948 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 VGND 0.030153f
C1949 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 VGND 0.234486f
C1950 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n16 VGND 0.050613f
C1951 tdc_0.vernier_delay_line_0.start_neg.t7 VGND 0.153672f
C1952 tdc_0.vernier_delay_line_0.start_neg.t6 VGND 0.047491f
C1953 tdc_0.vernier_delay_line_0.start_neg.n0 VGND 0.42006f
C1954 tdc_0.vernier_delay_line_0.start_neg.t8 VGND 0.061832f
C1955 tdc_0.vernier_delay_line_0.start_neg.t15 VGND 0.019725f
C1956 tdc_0.vernier_delay_line_0.start_neg.n1 VGND 0.043367f
C1957 tdc_0.vernier_delay_line_0.start_neg.t14 VGND 0.061832f
C1958 tdc_0.vernier_delay_line_0.start_neg.t13 VGND 0.019725f
C1959 tdc_0.vernier_delay_line_0.start_neg.n2 VGND 0.043087f
C1960 tdc_0.vernier_delay_line_0.start_neg.n3 VGND 0.013896f
C1961 tdc_0.vernier_delay_line_0.start_neg.t12 VGND 0.061832f
C1962 tdc_0.vernier_delay_line_0.start_neg.t10 VGND 0.019725f
C1963 tdc_0.vernier_delay_line_0.start_neg.n4 VGND 0.043367f
C1964 tdc_0.vernier_delay_line_0.start_neg.t11 VGND 0.061832f
C1965 tdc_0.vernier_delay_line_0.start_neg.t9 VGND 0.019725f
C1966 tdc_0.vernier_delay_line_0.start_neg.n5 VGND 0.043087f
C1967 tdc_0.vernier_delay_line_0.start_neg.n6 VGND 0.013747f
C1968 tdc_0.vernier_delay_line_0.start_neg.n7 VGND 0.187263f
C1969 tdc_0.vernier_delay_line_0.start_neg.t3 VGND 0.040569f
C1970 tdc_0.vernier_delay_line_0.start_neg.t4 VGND 0.040569f
C1971 tdc_0.vernier_delay_line_0.start_neg.n8 VGND 0.086755f
C1972 tdc_0.vernier_delay_line_0.start_neg.t1 VGND 0.013523f
C1973 tdc_0.vernier_delay_line_0.start_neg.t2 VGND 0.013523f
C1974 tdc_0.vernier_delay_line_0.start_neg.n9 VGND 0.029358f
C1975 tdc_0.vernier_delay_line_0.start_neg.n10 VGND 0.348878f
C1976 tdc_0.vernier_delay_line_0.start_neg.t5 VGND 0.153672f
C1977 tdc_0.vernier_delay_line_0.start_neg.t0 VGND 0.047491f
C1978 tdc_0.vernier_delay_line_0.start_neg.n11 VGND 0.369312f
C1979 tdc_0.vernier_delay_line_0.start_neg.n12 VGND 0.079715f
C1980 uio_in[0].t1 VGND 0.072685f
C1981 uio_in[0].t5 VGND 0.078634f
C1982 uio_in[0].n0 VGND 0.077149f
C1983 uio_in[0].t7 VGND 0.078369f
C1984 uio_in[0].n1 VGND 0.053689f
C1985 uio_in[0].t0 VGND 0.022787f
C1986 uio_in[0].t2 VGND 0.029248f
C1987 uio_in[0].t6 VGND 0.029248f
C1988 uio_in[0].n2 VGND 0.087662f
C1989 uio_in[0].n3 VGND 0.531341f
C1990 uio_in[0].n4 VGND 5.469f
C1991 uio_in[0].t3 VGND 0.073684f
C1992 uio_in[0].t4 VGND 0.023785f
C1993 uio_in[0].n5 VGND 0.074548f
C1994 uio_in[0].n6 VGND 0.62346f
C1995 ui_in[6].t0 VGND 0.064986f
C1996 ui_in[6].t1 VGND 0.070305f
C1997 ui_in[6].n0 VGND 0.068977f
C1998 ui_in[6].t5 VGND 0.070068f
C1999 ui_in[6].n1 VGND 0.048001f
C2000 ui_in[6].t6 VGND 0.020373f
C2001 ui_in[6].t7 VGND 0.02615f
C2002 ui_in[6].t4 VGND 0.02615f
C2003 ui_in[6].n2 VGND 0.078377f
C2004 ui_in[6].n3 VGND 0.397332f
C2005 ui_in[6].n4 VGND 4.07223f
C2006 ui_in[6].t2 VGND 0.065879f
C2007 ui_in[6].t3 VGND 0.021265f
C2008 ui_in[6].n5 VGND 0.066651f
C2009 ui_in[6].n6 VGND 0.565747f
C2010 ui_in[7].t1 VGND 0.08368f
C2011 ui_in[7].t5 VGND 0.090529f
C2012 ui_in[7].n0 VGND 0.088818f
C2013 ui_in[7].t7 VGND 0.090223f
C2014 ui_in[7].n1 VGND 0.06181f
C2015 ui_in[7].t0 VGND 0.026234f
C2016 ui_in[7].t4 VGND 0.033672f
C2017 ui_in[7].t6 VGND 0.033672f
C2018 ui_in[7].n2 VGND 0.100922f
C2019 ui_in[7].n3 VGND 0.609031f
C2020 ui_in[7].n4 VGND 5.81591f
C2021 ui_in[7].t2 VGND 0.084829f
C2022 ui_in[7].t3 VGND 0.027383f
C2023 ui_in[7].n5 VGND 0.085824f
C2024 ui_in[7].n6 VGND 0.719999f
C2025 tdc_0.vernier_delay_line_0.start_pos.t11 VGND 0.086445f
C2026 tdc_0.vernier_delay_line_0.start_pos.t9 VGND 0.027576f
C2027 tdc_0.vernier_delay_line_0.start_pos.n0 VGND 0.060238f
C2028 tdc_0.vernier_delay_line_0.start_pos.t8 VGND 0.086445f
C2029 tdc_0.vernier_delay_line_0.start_pos.t15 VGND 0.027576f
C2030 tdc_0.vernier_delay_line_0.start_pos.n1 VGND 0.060629f
C2031 tdc_0.vernier_delay_line_0.start_pos.n2 VGND 0.01943f
C2032 tdc_0.vernier_delay_line_0.start_pos.t14 VGND 0.086445f
C2033 tdc_0.vernier_delay_line_0.start_pos.t13 VGND 0.027576f
C2034 tdc_0.vernier_delay_line_0.start_pos.n3 VGND 0.060629f
C2035 tdc_0.vernier_delay_line_0.start_pos.t12 VGND 0.086445f
C2036 tdc_0.vernier_delay_line_0.start_pos.t10 VGND 0.027576f
C2037 tdc_0.vernier_delay_line_0.start_pos.n4 VGND 0.060238f
C2038 tdc_0.vernier_delay_line_0.start_pos.n5 VGND 0.019219f
C2039 tdc_0.vernier_delay_line_0.start_pos.n6 VGND 0.507295f
C2040 tdc_0.vernier_delay_line_0.start_pos.t0 VGND 0.069183f
C2041 tdc_0.vernier_delay_line_0.start_pos.t1 VGND 0.209408f
C2042 tdc_0.vernier_delay_line_0.start_pos.n7 VGND 0.531486f
C2043 tdc_0.vernier_delay_line_0.start_pos.n8 VGND 0.276923f
C2044 tdc_0.vernier_delay_line_0.start_pos.t3 VGND 0.018906f
C2045 tdc_0.vernier_delay_line_0.start_pos.t4 VGND 0.018906f
C2046 tdc_0.vernier_delay_line_0.start_pos.n9 VGND 0.044282f
C2047 tdc_0.vernier_delay_line_0.start_pos.t5 VGND 0.056718f
C2048 tdc_0.vernier_delay_line_0.start_pos.t6 VGND 0.056718f
C2049 tdc_0.vernier_delay_line_0.start_pos.n10 VGND 0.115544f
C2050 tdc_0.vernier_delay_line_0.start_pos.n11 VGND 0.480734f
C2051 tdc_0.vernier_delay_line_0.start_pos.t2 VGND 0.069203f
C2052 tdc_0.vernier_delay_line_0.start_pos.t7 VGND 0.209408f
C2053 tdc_0.vernier_delay_line_0.start_pos.n12 VGND 0.51072f
C2054 tdc_0.vernier_delay_line_0.start_pos.n13 VGND 0.261208f
C2055 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t1 VGND 0.165681f
C2056 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t0 VGND 0.051203f
C2057 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n0 VGND 0.451103f
C2058 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t8 VGND 0.066664f
C2059 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t14 VGND 0.021266f
C2060 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n1 VGND 0.046756f
C2061 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t13 VGND 0.066664f
C2062 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t11 VGND 0.021266f
C2063 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n2 VGND 0.046454f
C2064 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n3 VGND 0.014982f
C2065 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t12 VGND 0.066664f
C2066 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t10 VGND 0.021266f
C2067 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n4 VGND 0.046756f
C2068 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t9 VGND 0.066664f
C2069 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t15 VGND 0.021266f
C2070 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n5 VGND 0.046454f
C2071 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n6 VGND 0.014821f
C2072 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n7 VGND 0.229513f
C2073 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t7 VGND 0.043739f
C2074 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t5 VGND 0.043739f
C2075 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n8 VGND 0.093535f
C2076 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t2 VGND 0.01458f
C2077 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t3 VGND 0.01458f
C2078 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n9 VGND 0.031652f
C2079 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n10 VGND 0.376142f
C2080 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t6 VGND 0.165681f
C2081 tdc_0.diff_gen_0.delay_unit_2_6.in_2.t4 VGND 0.051203f
C2082 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n11 VGND 0.398173f
C2083 tdc_0.diff_gen_0.delay_unit_2_6.in_2.n12 VGND 0.085944f
C2084 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 VGND 0.059856f
C2085 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 VGND 0.019094f
C2086 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2087 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 VGND 0.059856f
C2088 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 VGND 0.019094f
C2089 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2090 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2091 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 VGND 0.059856f
C2092 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 VGND 0.019094f
C2093 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2094 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 VGND 0.059856f
C2095 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 VGND 0.019094f
C2096 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2097 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2098 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2099 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 VGND 0.047903f
C2100 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 VGND 0.144997f
C2101 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2102 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 VGND 0.191745f
C2103 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 VGND 0.013091f
C2104 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 VGND 0.013091f
C2105 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 VGND 0.030662f
C2106 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 VGND 0.039272f
C2107 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 VGND 0.039272f
C2108 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 VGND 0.080004f
C2109 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 VGND 0.332866f
C2110 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 VGND 0.060722f
C2111 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 VGND 0.060722f
C2112 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 VGND 0.070899f
C2113 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 VGND 0.060722f
C2114 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 VGND 0.060722f
C2115 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 VGND 0.070523f
C2116 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 VGND 0.632153f
C2117 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 VGND 0.045973f
C2118 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 VGND 0.156775f
C2119 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 VGND 0.144997f
C2120 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 VGND 0.240639f
C2121 tdc_0.vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 VGND 0.180864f
C2122 ui_in[4].t3 VGND 0.039584f
C2123 ui_in[4].t5 VGND 0.012778f
C2124 ui_in[4].n0 VGND 0.040049f
C2125 ui_in[4].t0 VGND 0.039048f
C2126 ui_in[4].t2 VGND 0.042244f
C2127 ui_in[4].n1 VGND 0.041446f
C2128 ui_in[4].t6 VGND 0.042102f
C2129 ui_in[4].n2 VGND 0.028843f
C2130 ui_in[4].t7 VGND 0.012242f
C2131 ui_in[4].t1 VGND 0.015712f
C2132 ui_in[4].t4 VGND 0.015712f
C2133 ui_in[4].n3 VGND 0.047094f
C2134 ui_in[4].n4 VGND 0.28086f
C2135 ui_in[4].n5 VGND 1.95509f
C2136 ui_in[4].n6 VGND 0.343484f
C2137 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 VGND 0.059856f
C2138 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 VGND 0.019094f
C2139 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2140 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 VGND 0.059856f
C2141 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 VGND 0.019094f
C2142 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2143 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2144 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 VGND 0.059856f
C2145 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 VGND 0.019094f
C2146 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2147 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 VGND 0.059856f
C2148 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 VGND 0.019094f
C2149 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2150 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2151 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2152 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 VGND 0.047903f
C2153 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 VGND 0.144997f
C2154 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2155 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 VGND 0.013091f
C2156 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 VGND 0.013091f
C2157 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 VGND 0.030662f
C2158 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 VGND 0.039272f
C2159 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 VGND 0.039272f
C2160 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 VGND 0.080004f
C2161 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 VGND 0.332866f
C2162 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 VGND 0.060722f
C2163 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 VGND 0.060722f
C2164 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 VGND 0.070899f
C2165 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 VGND 0.060722f
C2166 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 VGND 0.060722f
C2167 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 VGND 0.070523f
C2168 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 VGND 0.632153f
C2169 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 VGND 0.045973f
C2170 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 VGND 0.156775f
C2171 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 VGND 0.144997f
C2172 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 VGND 0.240639f
C2173 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 VGND 0.180864f
C2174 variable_delay_short_0.variable_delay_unit_4.in.t4 VGND 0.017058f
C2175 variable_delay_short_0.variable_delay_unit_4.in.t5 VGND 0.044984f
C2176 variable_delay_short_0.variable_delay_unit_4.in.n0 VGND 0.04731f
C2177 variable_delay_short_0.variable_delay_unit_4.in.t0 VGND 0.033139f
C2178 variable_delay_short_0.variable_delay_unit_4.in.t1 VGND 0.105354f
C2179 variable_delay_short_0.variable_delay_unit_4.in.n1 VGND 0.255341f
C2180 variable_delay_short_0.variable_delay_unit_4.in.t2 VGND 0.042943f
C2181 variable_delay_short_0.variable_delay_unit_4.in.t3 VGND 0.013862f
C2182 variable_delay_short_0.variable_delay_unit_4.in.n2 VGND 0.045161f
C2183 variable_delay_short_0.variable_delay_unit_4.in.n3 VGND 0.418008f
C2184 variable_delay_short_0.variable_delay_unit_3.in.t4 VGND 0.017058f
C2185 variable_delay_short_0.variable_delay_unit_3.in.t5 VGND 0.044984f
C2186 variable_delay_short_0.variable_delay_unit_3.in.n0 VGND 0.04731f
C2187 variable_delay_short_0.variable_delay_unit_3.in.t0 VGND 0.033139f
C2188 variable_delay_short_0.variable_delay_unit_3.in.t1 VGND 0.105354f
C2189 variable_delay_short_0.variable_delay_unit_3.in.n1 VGND 0.255341f
C2190 variable_delay_short_0.variable_delay_unit_3.in.t2 VGND 0.042943f
C2191 variable_delay_short_0.variable_delay_unit_3.in.t3 VGND 0.013862f
C2192 variable_delay_short_0.variable_delay_unit_3.in.n2 VGND 0.045161f
C2193 variable_delay_short_0.variable_delay_unit_3.in.n3 VGND 0.418008f
C2194 a_10108_23980.t1 VGND 0.059028f
C2195 a_10108_23980.t0 VGND 0.059028f
C2196 a_10108_23980.t2 VGND 0.059028f
C2197 a_10108_23980.n0 VGND 0.136068f
C2198 a_10108_23980.t4 VGND 0.059028f
C2199 a_10108_23980.t5 VGND 0.059028f
C2200 a_10108_23980.n1 VGND 0.139449f
C2201 a_10108_23980.n2 VGND 1.11221f
C2202 a_10108_23980.n3 VGND 0.258102f
C2203 a_10108_23980.t3 VGND 0.059028f
C2204 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 VGND 0.025758f
C2205 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 VGND 0.025758f
C2206 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 VGND 0.055083f
C2207 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 VGND 0.008586f
C2208 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 VGND 0.008586f
C2209 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 VGND 0.01864f
C2210 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 VGND 0.221512f
C2211 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 VGND 0.09757f
C2212 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 VGND 0.030153f
C2213 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 VGND 0.234486f
C2214 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 VGND 0.046129f
C2215 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 VGND 0.046129f
C2216 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 VGND 0.054044f
C2217 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 VGND 0.046129f
C2218 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 VGND 0.046129f
C2219 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 VGND 0.0538f
C2220 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 VGND 0.495704f
C2221 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 VGND 0.09757f
C2222 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 VGND 0.030153f
C2223 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 VGND 0.265657f
C2224 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 VGND 0.039259f
C2225 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 VGND 0.012524f
C2226 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 VGND 0.027534f
C2227 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 VGND 0.039259f
C2228 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 VGND 0.012524f
C2229 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 VGND 0.027357f
C2230 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 VGND 0.008823f
C2231 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 VGND 0.039259f
C2232 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2233 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 VGND 0.027534f
C2234 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2235 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 VGND 0.012524f
C2236 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 VGND 0.027357f
C2237 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 VGND 0.008728f
C2238 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 VGND 0.135162f
C2239 a_10958_30210.t3 VGND 0.024913f
C2240 a_10958_30210.t0 VGND 0.024913f
C2241 a_10958_30210.t2 VGND 0.024913f
C2242 a_10958_30210.n0 VGND 0.059872f
C2243 a_10958_30210.t12 VGND 0.096748f
C2244 a_10958_30210.t5 VGND 0.024913f
C2245 a_10958_30210.t9 VGND 0.024913f
C2246 a_10958_30210.n1 VGND 0.060504f
C2247 a_10958_30210.n2 VGND 0.369187f
C2248 a_10958_30210.t11 VGND 0.024913f
C2249 a_10958_30210.t7 VGND 0.024913f
C2250 a_10958_30210.n3 VGND 0.060504f
C2251 a_10958_30210.n4 VGND 0.182084f
C2252 a_10958_30210.t8 VGND 0.024913f
C2253 a_10958_30210.t10 VGND 0.024913f
C2254 a_10958_30210.n5 VGND 0.060504f
C2255 a_10958_30210.n6 VGND 0.221492f
C2256 a_10958_30210.t1 VGND 0.024913f
C2257 a_10958_30210.t6 VGND 0.024913f
C2258 a_10958_30210.n7 VGND 0.052659f
C2259 a_10958_30210.n8 VGND 0.137512f
C2260 a_10958_30210.n9 VGND 0.342225f
C2261 a_10958_30210.n10 VGND 0.057757f
C2262 a_10958_30210.t4 VGND 0.024913f
C2263 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 VGND 0.059856f
C2264 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 VGND 0.019094f
C2265 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2266 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 VGND 0.059856f
C2267 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 VGND 0.019094f
C2268 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2269 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2270 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 VGND 0.059856f
C2271 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 VGND 0.019094f
C2272 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2273 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 VGND 0.059856f
C2274 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 VGND 0.019094f
C2275 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2276 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2277 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2278 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 VGND 0.047903f
C2279 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 VGND 0.144997f
C2280 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2281 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 VGND 0.013091f
C2282 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 VGND 0.013091f
C2283 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 VGND 0.030662f
C2284 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 VGND 0.039272f
C2285 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 VGND 0.039272f
C2286 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 VGND 0.080004f
C2287 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 VGND 0.332866f
C2288 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 VGND 0.060722f
C2289 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 VGND 0.060722f
C2290 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 VGND 0.070899f
C2291 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 VGND 0.060722f
C2292 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 VGND 0.060722f
C2293 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 VGND 0.070523f
C2294 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 VGND 0.632153f
C2295 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 VGND 0.045973f
C2296 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 VGND 0.156775f
C2297 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 VGND 0.144997f
C2298 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 VGND 0.240639f
C2299 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 VGND 0.180864f
C2300 variable_delay_short_0.variable_delay_unit_5.forward.t2 VGND 0.025654f
C2301 variable_delay_short_0.variable_delay_unit_5.forward.t3 VGND 0.067654f
C2302 variable_delay_short_0.variable_delay_unit_5.forward.n0 VGND 0.071153f
C2303 variable_delay_short_0.variable_delay_unit_5.forward.t0 VGND 0.04984f
C2304 variable_delay_short_0.variable_delay_unit_5.forward.t1 VGND 0.15845f
C2305 variable_delay_short_0.variable_delay_unit_5.forward.n1 VGND 0.384027f
C2306 variable_delay_short_0.variable_delay_unit_5.forward.n2 VGND 0.628675f
C2307 variable_delay_short_0.variable_delay_unit_5.in.t4 VGND 0.021119f
C2308 variable_delay_short_0.variable_delay_unit_5.in.t5 VGND 0.055694f
C2309 variable_delay_short_0.variable_delay_unit_5.in.n0 VGND 0.058574f
C2310 variable_delay_short_0.variable_delay_unit_5.in.t1 VGND 0.041029f
C2311 variable_delay_short_0.variable_delay_unit_5.in.t0 VGND 0.130438f
C2312 variable_delay_short_0.variable_delay_unit_5.in.n1 VGND 0.316137f
C2313 variable_delay_short_0.variable_delay_unit_5.in.t2 VGND 0.053167f
C2314 variable_delay_short_0.variable_delay_unit_5.in.t3 VGND 0.017162f
C2315 variable_delay_short_0.variable_delay_unit_5.in.n2 VGND 0.055913f
C2316 variable_delay_short_0.variable_delay_unit_5.in.n3 VGND 0.517534f
C2317 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C2318 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C2319 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.087567f
C2320 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.039734f
C2321 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C2322 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.202442f
C2323 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C2324 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.054262f
C2325 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.115417f
C2326 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.089004f
C2327 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C2328 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C2329 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.041221f
C2330 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.095888f
C2331 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C2332 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.108461f
C2333 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C2334 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 VGND 0.09757f
C2335 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 VGND 0.030153f
C2336 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2337 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 VGND 0.039259f
C2338 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 VGND 0.012524f
C2339 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2340 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 VGND 0.039259f
C2341 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 VGND 0.012524f
C2342 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2343 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2344 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 VGND 0.039259f
C2345 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2346 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2347 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2348 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 VGND 0.012524f
C2349 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2350 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2351 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2352 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 VGND 0.046129f
C2353 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 VGND 0.046129f
C2354 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2355 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 VGND 0.046129f
C2356 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2357 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2358 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2359 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 VGND 0.025758f
C2360 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 VGND 0.025758f
C2361 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2362 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 VGND 0.008586f
C2363 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 VGND 0.008586f
C2364 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2365 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2366 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 VGND 0.09757f
C2367 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 VGND 0.030153f
C2368 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2369 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t9 VGND 0.086195f
C2370 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t15 VGND 0.027496f
C2371 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n0 VGND 0.060063f
C2372 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t13 VGND 0.086195f
C2373 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t12 VGND 0.027496f
C2374 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n1 VGND 0.060453f
C2375 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n2 VGND 0.019374f
C2376 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t11 VGND 0.086195f
C2377 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t10 VGND 0.027496f
C2378 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n3 VGND 0.060453f
C2379 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t8 VGND 0.086195f
C2380 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t14 VGND 0.027496f
C2381 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n4 VGND 0.060063f
C2382 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n5 VGND 0.019163f
C2383 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n6 VGND 0.505822f
C2384 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t6 VGND 0.068982f
C2385 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t7 VGND 0.2088f
C2386 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n7 VGND 0.529943f
C2387 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n8 VGND 0.27612f
C2388 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t1 VGND 0.018851f
C2389 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t2 VGND 0.018851f
C2390 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n9 VGND 0.044154f
C2391 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t3 VGND 0.056553f
C2392 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t4 VGND 0.056553f
C2393 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n10 VGND 0.115209f
C2394 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n11 VGND 0.479339f
C2395 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t0 VGND 0.069002f
C2396 tdc_0.diff_gen_0.delay_unit_2_1.in_1.t5 VGND 0.2088f
C2397 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n12 VGND 0.509237f
C2398 tdc_0.diff_gen_0.delay_unit_2_1.in_1.n13 VGND 0.26045f
C2399 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 VGND 0.061913f
C2400 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 VGND 0.061913f
C2401 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 VGND 0.072289f
C2402 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 VGND 0.061913f
C2403 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 VGND 0.061913f
C2404 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 VGND 0.071905f
C2405 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 VGND 0.644548f
C2406 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 VGND 0.061029f
C2407 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 VGND 0.019469f
C2408 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 VGND 0.042527f
C2409 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 VGND 0.061029f
C2410 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 VGND 0.019469f
C2411 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 VGND 0.042803f
C2412 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 VGND 0.013718f
C2413 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 VGND 0.061029f
C2414 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 VGND 0.019469f
C2415 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 VGND 0.042803f
C2416 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 VGND 0.061029f
C2417 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 VGND 0.019469f
C2418 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 VGND 0.042527f
C2419 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 VGND 0.013568f
C2420 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 VGND 0.358144f
C2421 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 VGND 0.048842f
C2422 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 VGND 0.14784f
C2423 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 VGND 0.375222f
C2424 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 VGND 0.013347f
C2425 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 VGND 0.013347f
C2426 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 VGND 0.031263f
C2427 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 VGND 0.040042f
C2428 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 VGND 0.040042f
C2429 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 VGND 0.081573f
C2430 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 VGND 0.339393f
C2431 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 VGND 0.18441f
C2432 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 VGND 0.14784f
C2433 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 VGND 0.245357f
C2434 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 VGND 0.046875f
C2435 tdc_0.vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 VGND 0.159849f
C2436 a_10958_32492.t7 VGND 0.024913f
C2437 a_10958_32492.t5 VGND 0.096748f
C2438 a_10958_32492.t4 VGND 0.024913f
C2439 a_10958_32492.t6 VGND 0.024913f
C2440 a_10958_32492.n0 VGND 0.060504f
C2441 a_10958_32492.n1 VGND 0.369187f
C2442 a_10958_32492.t0 VGND 0.024913f
C2443 a_10958_32492.t3 VGND 0.024913f
C2444 a_10958_32492.n2 VGND 0.060504f
C2445 a_10958_32492.n3 VGND 0.182084f
C2446 a_10958_32492.t2 VGND 0.024913f
C2447 a_10958_32492.t1 VGND 0.024913f
C2448 a_10958_32492.n4 VGND 0.060504f
C2449 a_10958_32492.n5 VGND 0.221492f
C2450 a_10958_32492.t10 VGND 0.024913f
C2451 a_10958_32492.t12 VGND 0.024913f
C2452 a_10958_32492.n6 VGND 0.052659f
C2453 a_10958_32492.n7 VGND 0.137512f
C2454 a_10958_32492.t8 VGND 0.024913f
C2455 a_10958_32492.t9 VGND 0.024913f
C2456 a_10958_32492.n8 VGND 0.057757f
C2457 a_10958_32492.n9 VGND 0.342225f
C2458 a_10958_32492.n10 VGND 0.059872f
C2459 a_10958_32492.t11 VGND 0.024913f
C2460 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t11 VGND 0.086195f
C2461 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t9 VGND 0.027496f
C2462 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n0 VGND 0.060063f
C2463 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t8 VGND 0.086195f
C2464 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t15 VGND 0.027496f
C2465 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n1 VGND 0.060453f
C2466 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n2 VGND 0.019374f
C2467 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t14 VGND 0.086195f
C2468 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t13 VGND 0.027496f
C2469 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n3 VGND 0.060453f
C2470 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t12 VGND 0.086195f
C2471 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t10 VGND 0.027496f
C2472 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n4 VGND 0.060063f
C2473 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n5 VGND 0.019163f
C2474 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n6 VGND 0.505822f
C2475 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t6 VGND 0.068982f
C2476 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t7 VGND 0.2088f
C2477 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n7 VGND 0.529943f
C2478 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n8 VGND 0.27612f
C2479 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t2 VGND 0.018851f
C2480 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t0 VGND 0.018851f
C2481 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n9 VGND 0.044154f
C2482 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t4 VGND 0.056553f
C2483 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t5 VGND 0.056553f
C2484 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n10 VGND 0.115209f
C2485 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n11 VGND 0.479339f
C2486 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t1 VGND 0.069002f
C2487 tdc_0.diff_gen_0.delay_unit_2_3.in_1.t3 VGND 0.2088f
C2488 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n12 VGND 0.509237f
C2489 tdc_0.diff_gen_0.delay_unit_2_3.in_1.n13 VGND 0.26045f
C2490 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t3 VGND 0.165681f
C2491 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t2 VGND 0.051203f
C2492 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n0 VGND 0.451103f
C2493 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t13 VGND 0.066664f
C2494 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t11 VGND 0.021266f
C2495 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n1 VGND 0.046756f
C2496 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t10 VGND 0.066664f
C2497 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t8 VGND 0.021266f
C2498 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n2 VGND 0.046454f
C2499 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n3 VGND 0.014982f
C2500 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t9 VGND 0.066664f
C2501 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t15 VGND 0.021266f
C2502 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n4 VGND 0.046756f
C2503 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t14 VGND 0.066664f
C2504 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t12 VGND 0.021266f
C2505 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n5 VGND 0.046454f
C2506 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n6 VGND 0.014821f
C2507 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n7 VGND 0.229513f
C2508 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t4 VGND 0.043739f
C2509 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t5 VGND 0.043739f
C2510 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n8 VGND 0.093535f
C2511 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t0 VGND 0.01458f
C2512 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t6 VGND 0.01458f
C2513 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n9 VGND 0.031652f
C2514 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n10 VGND 0.376142f
C2515 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t1 VGND 0.165681f
C2516 tdc_0.diff_gen_0.delay_unit_2_2.in_2.t7 VGND 0.051203f
C2517 tdc_0.diff_gen_0.delay_unit_2_2.in_2.n11 VGND 0.398173f
C2518 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t4 VGND 0.027086f
C2519 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t6 VGND 0.034765f
C2520 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t2 VGND 0.034765f
C2521 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n0 VGND 0.10415f
C2522 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t0 VGND 0.067642f
C2523 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t1 VGND 0.215011f
C2524 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n1 VGND 0.85898f
C2525 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t5 VGND 0.093153f
C2526 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t3 VGND 0.086397f
C2527 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.t7 VGND 0.093468f
C2528 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n2 VGND 0.091702f
C2529 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n3 VGND 0.063806f
C2530 variable_delay_dummy_0.variable_delay_unit_0.tristate_inverter_1.en.n4 VGND 0.942937f
C2531 uo_out[3].t5 VGND 0.007815f
C2532 uo_out[3].t4 VGND 0.026417f
C2533 uo_out[3].n0 VGND 0.021415f
C2534 uo_out[3].t0 VGND 0.015221f
C2535 uo_out[3].t3 VGND 0.015221f
C2536 uo_out[3].n1 VGND 0.032348f
C2537 uo_out[3].n2 VGND 0.141125f
C2538 uo_out[3].t2 VGND 0.005074f
C2539 uo_out[3].t1 VGND 0.005074f
C2540 uo_out[3].n3 VGND 0.011015f
C2541 uo_out[3].n4 VGND 0.037476f
C2542 uo_out[3].n5 VGND 0.713178f
C2543 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 VGND 0.930597f
C2544 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.400887f
C2545 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 VGND 1.11317f
C2546 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.087567f
C2547 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C2548 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.097942f
C2549 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.089004f
C2550 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.08317f
C2551 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C2552 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.041221f
C2553 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.095888f
C2554 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C2555 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.108461f
C2556 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C2557 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C2558 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C2559 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 VGND 0.115417f
C2560 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C2561 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C2562 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.041341f
C2563 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.096169f
C2564 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C2565 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.089265f
C2566 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.083414f
C2567 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C2568 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.202074f
C2569 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.087824f
C2570 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.03985f
C2571 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C2572 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.200787f
C2573 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C2574 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.054421f
C2575 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C2576 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C2577 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.107523f
C2578 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C2579 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C2580 a_10958_25646.t10 VGND 0.024913f
C2581 a_10958_25646.t5 VGND 0.096748f
C2582 a_10958_25646.t2 VGND 0.024913f
C2583 a_10958_25646.t6 VGND 0.024913f
C2584 a_10958_25646.n0 VGND 0.060504f
C2585 a_10958_25646.n1 VGND 0.369187f
C2586 a_10958_25646.t4 VGND 0.024913f
C2587 a_10958_25646.t1 VGND 0.024913f
C2588 a_10958_25646.n2 VGND 0.060504f
C2589 a_10958_25646.n3 VGND 0.182084f
C2590 a_10958_25646.t0 VGND 0.024913f
C2591 a_10958_25646.t7 VGND 0.024913f
C2592 a_10958_25646.n4 VGND 0.060504f
C2593 a_10958_25646.n5 VGND 0.221492f
C2594 a_10958_25646.t12 VGND 0.024913f
C2595 a_10958_25646.t3 VGND 0.024913f
C2596 a_10958_25646.n6 VGND 0.052659f
C2597 a_10958_25646.n7 VGND 0.137512f
C2598 a_10958_25646.t8 VGND 0.024913f
C2599 a_10958_25646.t9 VGND 0.024913f
C2600 a_10958_25646.n8 VGND 0.057757f
C2601 a_10958_25646.n9 VGND 0.342225f
C2602 a_10958_25646.n10 VGND 0.059872f
C2603 a_10958_25646.t11 VGND 0.024913f
C2604 uo_out[0].t4 VGND 0.007317f
C2605 uo_out[0].t5 VGND 0.024735f
C2606 uo_out[0].n0 VGND 0.020051f
C2607 uo_out[0].t1 VGND 0.014251f
C2608 uo_out[0].t3 VGND 0.014251f
C2609 uo_out[0].n1 VGND 0.030287f
C2610 uo_out[0].n2 VGND 0.132137f
C2611 uo_out[0].t2 VGND 0.004751f
C2612 uo_out[0].t0 VGND 0.004751f
C2613 uo_out[0].n3 VGND 0.010313f
C2614 uo_out[0].n4 VGND 0.03509f
C2615 uo_out[0].n5 VGND 1.00891f
C2616 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t8 VGND 0.086195f
C2617 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t14 VGND 0.027496f
C2618 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n0 VGND 0.060063f
C2619 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t13 VGND 0.086195f
C2620 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t12 VGND 0.027496f
C2621 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n1 VGND 0.060453f
C2622 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n2 VGND 0.019374f
C2623 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t11 VGND 0.086195f
C2624 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t10 VGND 0.027496f
C2625 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n3 VGND 0.060453f
C2626 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t9 VGND 0.086195f
C2627 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t15 VGND 0.027496f
C2628 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n4 VGND 0.060063f
C2629 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n5 VGND 0.019163f
C2630 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n6 VGND 0.505822f
C2631 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t0 VGND 0.068982f
C2632 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t1 VGND 0.2088f
C2633 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n7 VGND 0.529943f
C2634 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n8 VGND 0.27612f
C2635 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t3 VGND 0.018851f
C2636 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t4 VGND 0.018851f
C2637 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n9 VGND 0.044154f
C2638 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t6 VGND 0.056553f
C2639 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t7 VGND 0.056553f
C2640 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n10 VGND 0.115209f
C2641 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n11 VGND 0.479339f
C2642 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t2 VGND 0.069002f
C2643 tdc_0.diff_gen_0.delay_unit_2_6.in_1.t5 VGND 0.2088f
C2644 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n12 VGND 0.509237f
C2645 tdc_0.diff_gen_0.delay_unit_2_6.in_1.n13 VGND 0.26045f
C2646 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 VGND 0.09757f
C2647 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 VGND 0.030153f
C2648 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2649 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 VGND 0.039259f
C2650 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 VGND 0.012524f
C2651 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2652 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 VGND 0.039259f
C2653 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 VGND 0.012524f
C2654 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2655 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2656 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 VGND 0.039259f
C2657 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 VGND 0.012524f
C2658 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2659 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 VGND 0.039259f
C2660 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2661 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2662 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2663 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2664 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 VGND 0.046129f
C2665 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 VGND 0.046129f
C2666 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2667 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2668 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 VGND 0.046129f
C2669 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2670 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2671 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 VGND 0.025758f
C2672 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 VGND 0.025758f
C2673 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2674 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 VGND 0.008586f
C2675 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 VGND 0.008586f
C2676 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2677 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2678 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 VGND 0.09757f
C2679 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 VGND 0.030153f
C2680 tdc_0.vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2681 a_10108_30826.t0 VGND 0.059028f
C2682 a_10108_30826.t2 VGND 0.059028f
C2683 a_10108_30826.t5 VGND 0.059028f
C2684 a_10108_30826.n0 VGND 0.136068f
C2685 a_10108_30826.t3 VGND 0.059028f
C2686 a_10108_30826.t4 VGND 0.059028f
C2687 a_10108_30826.n1 VGND 0.258102f
C2688 a_10108_30826.n2 VGND 1.11221f
C2689 a_10108_30826.n3 VGND 0.139449f
C2690 a_10108_30826.t1 VGND 0.059028f
C2691 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 VGND 0.09757f
C2692 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 VGND 0.030153f
C2693 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2694 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 VGND 0.039259f
C2695 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 VGND 0.012524f
C2696 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2697 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 VGND 0.039259f
C2698 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 VGND 0.012524f
C2699 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2700 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2701 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2702 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 VGND 0.012524f
C2703 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2704 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 VGND 0.039259f
C2705 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 VGND 0.012524f
C2706 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2707 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2708 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2709 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 VGND 0.046129f
C2710 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 VGND 0.046129f
C2711 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2712 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2713 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 VGND 0.046129f
C2714 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2715 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2716 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 VGND 0.025758f
C2717 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 VGND 0.025758f
C2718 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2719 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 VGND 0.008586f
C2720 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 VGND 0.008586f
C2721 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2722 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2723 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 VGND 0.09757f
C2724 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 VGND 0.030153f
C2725 tdc_0.vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2726 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t4 VGND 0.027086f
C2727 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t5 VGND 0.034765f
C2728 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t7 VGND 0.034765f
C2729 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n0 VGND 0.10415f
C2730 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t0 VGND 0.067642f
C2731 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t1 VGND 0.215011f
C2732 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n1 VGND 0.85898f
C2733 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VGND 0.093153f
C2734 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t2 VGND 0.086397f
C2735 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VGND 0.093468f
C2736 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n2 VGND 0.091702f
C2737 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n3 VGND 0.063806f
C2738 variable_delay_dummy_0.variable_delay_unit_1.tristate_inverter_1.en.n4 VGND 0.942937f
C2739 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C2740 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C2741 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.087567f
C2742 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C2743 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C2744 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C2745 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C2746 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C2747 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.115417f
C2748 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.089004f
C2749 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C2750 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C2751 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.041221f
C2752 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.095888f
C2753 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C2754 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.108461f
C2755 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C2756 a_10958_27928.t5 VGND 0.024913f
C2757 a_10958_27928.t4 VGND 0.024913f
C2758 a_10958_27928.t7 VGND 0.024913f
C2759 a_10958_27928.n0 VGND 0.059872f
C2760 a_10958_27928.t12 VGND 0.096748f
C2761 a_10958_27928.t2 VGND 0.024913f
C2762 a_10958_27928.t9 VGND 0.024913f
C2763 a_10958_27928.n1 VGND 0.060504f
C2764 a_10958_27928.n2 VGND 0.369187f
C2765 a_10958_27928.t11 VGND 0.024913f
C2766 a_10958_27928.t0 VGND 0.024913f
C2767 a_10958_27928.n3 VGND 0.060504f
C2768 a_10958_27928.n4 VGND 0.182084f
C2769 a_10958_27928.t3 VGND 0.024913f
C2770 a_10958_27928.t10 VGND 0.024913f
C2771 a_10958_27928.n5 VGND 0.060504f
C2772 a_10958_27928.n6 VGND 0.221492f
C2773 a_10958_27928.t6 VGND 0.024913f
C2774 a_10958_27928.t1 VGND 0.024913f
C2775 a_10958_27928.n7 VGND 0.052659f
C2776 a_10958_27928.n8 VGND 0.137512f
C2777 a_10958_27928.n9 VGND 0.342225f
C2778 a_10958_27928.n10 VGND 0.057757f
C2779 a_10958_27928.t8 VGND 0.024913f
C2780 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t11 VGND 0.086195f
C2781 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t8 VGND 0.027496f
C2782 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n0 VGND 0.060063f
C2783 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t14 VGND 0.086195f
C2784 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t13 VGND 0.027496f
C2785 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n1 VGND 0.060453f
C2786 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n2 VGND 0.019374f
C2787 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t12 VGND 0.086195f
C2788 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t10 VGND 0.027496f
C2789 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n3 VGND 0.060453f
C2790 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t9 VGND 0.086195f
C2791 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t15 VGND 0.027496f
C2792 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n4 VGND 0.060063f
C2793 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n5 VGND 0.019163f
C2794 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n6 VGND 0.505822f
C2795 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t6 VGND 0.068982f
C2796 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t7 VGND 0.2088f
C2797 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n7 VGND 0.529943f
C2798 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n8 VGND 0.27612f
C2799 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t0 VGND 0.018851f
C2800 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t1 VGND 0.018851f
C2801 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n9 VGND 0.044154f
C2802 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t4 VGND 0.056553f
C2803 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t5 VGND 0.056553f
C2804 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n10 VGND 0.115209f
C2805 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n11 VGND 0.479339f
C2806 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t2 VGND 0.069002f
C2807 tdc_0.diff_gen_0.delay_unit_2_4.in_1.t3 VGND 0.2088f
C2808 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n12 VGND 0.509237f
C2809 tdc_0.diff_gen_0.delay_unit_2_4.in_1.n13 VGND 0.26045f
C2810 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t1 VGND 0.165681f
C2811 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t0 VGND 0.051203f
C2812 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n0 VGND 0.451103f
C2813 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t11 VGND 0.066664f
C2814 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t10 VGND 0.021266f
C2815 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n1 VGND 0.046756f
C2816 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t9 VGND 0.066664f
C2817 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t15 VGND 0.021266f
C2818 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n2 VGND 0.046454f
C2819 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n3 VGND 0.014982f
C2820 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t8 VGND 0.066664f
C2821 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t14 VGND 0.021266f
C2822 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n4 VGND 0.046756f
C2823 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t13 VGND 0.066664f
C2824 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t12 VGND 0.021266f
C2825 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n5 VGND 0.046454f
C2826 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n6 VGND 0.014821f
C2827 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n7 VGND 0.229513f
C2828 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t6 VGND 0.043739f
C2829 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t7 VGND 0.043739f
C2830 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n8 VGND 0.093535f
C2831 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t4 VGND 0.01458f
C2832 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t2 VGND 0.01458f
C2833 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n9 VGND 0.031652f
C2834 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n10 VGND 0.376142f
C2835 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t5 VGND 0.165681f
C2836 tdc_0.diff_gen_0.delay_unit_2_3.in_2.t3 VGND 0.051203f
C2837 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n11 VGND 0.398173f
C2838 tdc_0.diff_gen_0.delay_unit_2_3.in_2.n12 VGND 0.085944f
C2839 ui_in[5].t5 VGND 0.049226f
C2840 ui_in[5].t7 VGND 0.053255f
C2841 ui_in[5].n0 VGND 0.052248f
C2842 ui_in[5].t3 VGND 0.053075f
C2843 ui_in[5].n1 VGND 0.03636f
C2844 ui_in[5].t4 VGND 0.015432f
C2845 ui_in[5].t6 VGND 0.019808f
C2846 ui_in[5].t2 VGND 0.019808f
C2847 ui_in[5].n2 VGND 0.059369f
C2848 ui_in[5].n3 VGND 0.360373f
C2849 ui_in[5].n4 VGND 2.81694f
C2850 ui_in[5].t0 VGND 0.049902f
C2851 ui_in[5].t1 VGND 0.016108f
C2852 ui_in[5].n5 VGND 0.050487f
C2853 ui_in[5].n6 VGND 0.424074f
C2854 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t2 VGND 0.019446f
C2855 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t4 VGND 0.02496f
C2856 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t6 VGND 0.02496f
C2857 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n0 VGND 0.074774f
C2858 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t1 VGND 0.048564f
C2859 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t0 VGND 0.154367f
C2860 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n1 VGND 0.616703f
C2861 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t5 VGND 0.066879f
C2862 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t3 VGND 0.062029f
C2863 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.t7 VGND 0.067105f
C2864 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n2 VGND 0.065837f
C2865 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n3 VGND 0.045809f
C2866 variable_delay_short_0.variable_delay_unit_2.tristate_inverter_1.en.n4 VGND 0.676981f
C2867 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 VGND 0.059856f
C2868 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 VGND 0.019094f
C2869 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 VGND 0.041709f
C2870 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 VGND 0.059856f
C2871 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 VGND 0.019094f
C2872 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 VGND 0.04198f
C2873 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 VGND 0.013454f
C2874 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 VGND 0.059856f
C2875 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 VGND 0.019094f
C2876 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 VGND 0.04198f
C2877 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 VGND 0.059856f
C2878 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 VGND 0.019094f
C2879 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 VGND 0.041709f
C2880 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 VGND 0.013307f
C2881 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 VGND 0.351257f
C2882 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 VGND 0.047903f
C2883 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 VGND 0.144997f
C2884 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 VGND 0.368007f
C2885 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 VGND 0.191745f
C2886 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 VGND 0.013091f
C2887 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 VGND 0.013091f
C2888 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 VGND 0.030662f
C2889 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 VGND 0.039272f
C2890 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 VGND 0.039272f
C2891 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 VGND 0.080004f
C2892 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 VGND 0.332866f
C2893 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 VGND 0.060722f
C2894 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 VGND 0.060722f
C2895 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 VGND 0.070899f
C2896 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 VGND 0.060722f
C2897 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 VGND 0.060722f
C2898 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 VGND 0.070523f
C2899 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 VGND 0.632153f
C2900 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 VGND 0.045973f
C2901 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 VGND 0.156775f
C2902 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 VGND 0.144997f
C2903 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 VGND 0.240639f
C2904 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 VGND 0.180864f
C2905 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C2906 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.041341f
C2907 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.096169f
C2908 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C2909 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.089265f
C2910 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.083414f
C2911 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C2912 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.202074f
C2913 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.087824f
C2914 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C2915 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C2916 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.200787f
C2917 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.054421f
C2918 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C2919 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C2920 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C2921 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.107523f
C2922 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C2923 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C2924 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 VGND 0.09757f
C2925 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 VGND 0.030153f
C2926 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 VGND 0.265657f
C2927 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 VGND 0.039259f
C2928 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 VGND 0.012524f
C2929 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 VGND 0.027534f
C2930 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 VGND 0.039259f
C2931 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 VGND 0.012524f
C2932 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 VGND 0.027357f
C2933 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 VGND 0.008823f
C2934 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 VGND 0.039259f
C2935 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 VGND 0.012524f
C2936 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 VGND 0.027534f
C2937 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 VGND 0.039259f
C2938 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 VGND 0.012524f
C2939 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 VGND 0.027357f
C2940 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 VGND 0.008728f
C2941 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 VGND 0.135162f
C2942 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 VGND 0.046129f
C2943 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 VGND 0.046129f
C2944 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 VGND 0.054044f
C2945 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 VGND 0.046129f
C2946 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 VGND 0.046129f
C2947 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 VGND 0.0538f
C2948 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 VGND 0.495704f
C2949 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 VGND 0.025758f
C2950 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 VGND 0.025758f
C2951 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 VGND 0.055083f
C2952 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 VGND 0.008586f
C2953 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 VGND 0.008586f
C2954 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 VGND 0.01864f
C2955 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 VGND 0.221512f
C2956 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 VGND 0.09757f
C2957 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 VGND 0.030153f
C2958 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 VGND 0.234486f
C2959 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t7 VGND 0.165681f
C2960 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t6 VGND 0.051203f
C2961 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n0 VGND 0.451103f
C2962 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t8 VGND 0.066664f
C2963 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t15 VGND 0.021266f
C2964 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n1 VGND 0.046756f
C2965 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t14 VGND 0.066664f
C2966 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t12 VGND 0.021266f
C2967 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n2 VGND 0.046454f
C2968 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n3 VGND 0.014982f
C2969 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t13 VGND 0.066664f
C2970 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t11 VGND 0.021266f
C2971 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n4 VGND 0.046756f
C2972 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t10 VGND 0.066664f
C2973 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t9 VGND 0.021266f
C2974 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n5 VGND 0.046454f
C2975 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n6 VGND 0.014821f
C2976 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n7 VGND 0.229513f
C2977 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t4 VGND 0.043739f
C2978 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t2 VGND 0.043739f
C2979 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n8 VGND 0.093535f
C2980 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t1 VGND 0.01458f
C2981 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t3 VGND 0.01458f
C2982 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n9 VGND 0.031652f
C2983 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n10 VGND 0.376142f
C2984 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t5 VGND 0.165681f
C2985 tdc_0.diff_gen_0.delay_unit_2_4.in_2.t0 VGND 0.051203f
C2986 tdc_0.diff_gen_0.delay_unit_2_4.in_2.n11 VGND 0.398173f
C2987 a_10958_34774.t5 VGND 0.024913f
C2988 a_10958_34774.t6 VGND 0.024913f
C2989 a_10958_34774.t8 VGND 0.024913f
C2990 a_10958_34774.n0 VGND 0.059872f
C2991 a_10958_34774.t3 VGND 0.096748f
C2992 a_10958_34774.t12 VGND 0.024913f
C2993 a_10958_34774.t0 VGND 0.024913f
C2994 a_10958_34774.n1 VGND 0.060504f
C2995 a_10958_34774.n2 VGND 0.369187f
C2996 a_10958_34774.t2 VGND 0.024913f
C2997 a_10958_34774.t4 VGND 0.024913f
C2998 a_10958_34774.n3 VGND 0.060504f
C2999 a_10958_34774.n4 VGND 0.182084f
C3000 a_10958_34774.t10 VGND 0.024913f
C3001 a_10958_34774.t1 VGND 0.024913f
C3002 a_10958_34774.n5 VGND 0.060504f
C3003 a_10958_34774.n6 VGND 0.221492f
C3004 a_10958_34774.t7 VGND 0.024913f
C3005 a_10958_34774.t11 VGND 0.024913f
C3006 a_10958_34774.n7 VGND 0.052659f
C3007 a_10958_34774.n8 VGND 0.137512f
C3008 a_10958_34774.n9 VGND 0.342225f
C3009 a_10958_34774.n10 VGND 0.057757f
C3010 a_10958_34774.t9 VGND 0.024913f
C3011 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 VGND 0.060722f
C3012 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 VGND 0.060722f
C3013 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 VGND 0.070899f
C3014 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 VGND 0.060722f
C3015 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 VGND 0.060722f
C3016 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 VGND 0.070523f
C3017 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 VGND 0.632153f
C3018 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 VGND 0.059856f
C3019 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 VGND 0.019094f
C3020 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 VGND 0.041709f
C3021 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 VGND 0.059856f
C3022 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 VGND 0.019094f
C3023 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 VGND 0.04198f
C3024 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 VGND 0.013454f
C3025 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 VGND 0.059856f
C3026 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 VGND 0.019094f
C3027 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 VGND 0.04198f
C3028 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 VGND 0.059856f
C3029 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 VGND 0.019094f
C3030 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 VGND 0.041709f
C3031 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 VGND 0.013307f
C3032 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 VGND 0.351257f
C3033 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 VGND 0.047903f
C3034 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 VGND 0.144997f
C3035 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 VGND 0.368007f
C3036 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 VGND 0.013091f
C3037 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 VGND 0.013091f
C3038 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 VGND 0.030662f
C3039 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 VGND 0.039272f
C3040 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 VGND 0.039272f
C3041 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 VGND 0.080004f
C3042 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 VGND 0.332866f
C3043 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 VGND 0.180864f
C3044 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 VGND 0.144997f
C3045 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 VGND 0.240639f
C3046 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 VGND 0.045973f
C3047 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 VGND 0.156775f
C3048 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t12 VGND 0.086195f
C3049 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t10 VGND 0.027496f
C3050 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n0 VGND 0.060063f
C3051 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t9 VGND 0.086195f
C3052 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t15 VGND 0.027496f
C3053 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n1 VGND 0.060453f
C3054 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n2 VGND 0.019374f
C3055 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t14 VGND 0.086195f
C3056 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t13 VGND 0.027496f
C3057 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n3 VGND 0.060453f
C3058 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t11 VGND 0.086195f
C3059 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t8 VGND 0.027496f
C3060 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n4 VGND 0.060063f
C3061 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n5 VGND 0.019163f
C3062 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n6 VGND 0.505822f
C3063 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t0 VGND 0.068982f
C3064 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t1 VGND 0.2088f
C3065 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n7 VGND 0.529943f
C3066 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n8 VGND 0.302329f
C3067 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t5 VGND 0.018851f
C3068 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t2 VGND 0.018851f
C3069 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n9 VGND 0.044154f
C3070 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t3 VGND 0.056553f
C3071 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t6 VGND 0.056553f
C3072 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n10 VGND 0.115209f
C3073 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n11 VGND 0.479339f
C3074 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t4 VGND 0.069002f
C3075 tdc_0.diff_gen_0.delay_unit_2_5.in_1.t7 VGND 0.2088f
C3076 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n12 VGND 0.509237f
C3077 tdc_0.diff_gen_0.delay_unit_2_5.in_1.n13 VGND 0.26045f
C3078 tdc_0.diff_gen_0.delay_unit_2_4.out_1 VGND 0.212791f
C3079 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t2 VGND 0.165681f
C3080 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t3 VGND 0.051203f
C3081 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n0 VGND 0.451103f
C3082 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t14 VGND 0.066664f
C3083 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t13 VGND 0.021266f
C3084 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n1 VGND 0.046756f
C3085 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t12 VGND 0.066664f
C3086 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t10 VGND 0.021266f
C3087 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n2 VGND 0.046454f
C3088 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n3 VGND 0.014982f
C3089 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t11 VGND 0.066664f
C3090 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t9 VGND 0.021266f
C3091 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n4 VGND 0.046756f
C3092 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t8 VGND 0.066664f
C3093 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t15 VGND 0.021266f
C3094 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n5 VGND 0.046454f
C3095 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n6 VGND 0.014821f
C3096 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n7 VGND 0.229513f
C3097 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t4 VGND 0.043739f
C3098 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t0 VGND 0.043739f
C3099 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n8 VGND 0.093535f
C3100 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t1 VGND 0.01458f
C3101 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t5 VGND 0.01458f
C3102 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n9 VGND 0.031652f
C3103 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n10 VGND 0.376142f
C3104 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t6 VGND 0.165681f
C3105 tdc_0.diff_gen_0.delay_unit_2_5.in_2.t7 VGND 0.051203f
C3106 tdc_0.diff_gen_0.delay_unit_2_5.in_2.n11 VGND 0.398173f
C3107 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t13 VGND 0.086195f
C3108 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t11 VGND 0.027496f
C3109 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n0 VGND 0.060063f
C3110 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t10 VGND 0.086195f
C3111 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t9 VGND 0.027496f
C3112 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n1 VGND 0.060453f
C3113 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n2 VGND 0.019374f
C3114 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t8 VGND 0.086195f
C3115 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t15 VGND 0.027496f
C3116 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n3 VGND 0.060453f
C3117 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t14 VGND 0.086195f
C3118 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t12 VGND 0.027496f
C3119 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n4 VGND 0.060063f
C3120 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n5 VGND 0.019163f
C3121 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n6 VGND 0.505822f
C3122 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t0 VGND 0.068982f
C3123 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t1 VGND 0.2088f
C3124 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n7 VGND 0.529943f
C3125 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n8 VGND 0.27612f
C3126 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t3 VGND 0.018851f
C3127 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t4 VGND 0.018851f
C3128 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n9 VGND 0.044154f
C3129 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t5 VGND 0.056553f
C3130 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t6 VGND 0.056553f
C3131 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n10 VGND 0.115209f
C3132 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n11 VGND 0.479339f
C3133 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t2 VGND 0.069002f
C3134 tdc_0.diff_gen_0.delay_unit_2_2.in_1.t7 VGND 0.2088f
C3135 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n12 VGND 0.509237f
C3136 tdc_0.diff_gen_0.delay_unit_2_2.in_1.n13 VGND 0.26045f
C3137 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t0 VGND 0.165681f
C3138 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t7 VGND 0.051203f
C3139 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n0 VGND 0.451103f
C3140 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t8 VGND 0.066664f
C3141 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t14 VGND 0.021266f
C3142 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n1 VGND 0.046756f
C3143 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t13 VGND 0.066664f
C3144 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t11 VGND 0.021266f
C3145 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n2 VGND 0.046454f
C3146 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n3 VGND 0.014982f
C3147 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t12 VGND 0.066664f
C3148 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t10 VGND 0.021266f
C3149 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n4 VGND 0.046756f
C3150 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t9 VGND 0.066664f
C3151 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t15 VGND 0.021266f
C3152 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n5 VGND 0.046454f
C3153 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n6 VGND 0.014821f
C3154 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n7 VGND 0.229513f
C3155 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t6 VGND 0.043739f
C3156 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t4 VGND 0.043739f
C3157 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n8 VGND 0.093535f
C3158 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t1 VGND 0.01458f
C3159 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t2 VGND 0.01458f
C3160 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n9 VGND 0.031652f
C3161 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n10 VGND 0.376142f
C3162 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t5 VGND 0.165681f
C3163 tdc_0.diff_gen_0.delay_unit_2_1.in_2.t3 VGND 0.051203f
C3164 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n11 VGND 0.398173f
C3165 tdc_0.diff_gen_0.delay_unit_2_1.in_2.n12 VGND 0.085944f
C3166 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t2 VGND 0.019446f
C3167 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t4 VGND 0.02496f
C3168 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t6 VGND 0.02496f
C3169 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n0 VGND 0.074774f
C3170 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t1 VGND 0.048564f
C3171 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t0 VGND 0.154367f
C3172 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n1 VGND 0.616703f
C3173 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t5 VGND 0.066879f
C3174 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t3 VGND 0.062029f
C3175 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.t7 VGND 0.067105f
C3176 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n2 VGND 0.065837f
C3177 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n3 VGND 0.045809f
C3178 variable_delay_short_0.variable_delay_unit_4.tristate_inverter_1.en.n4 VGND 0.676981f
C3179 a_10108_26262.t5 VGND 0.059028f
C3180 a_10108_26262.t3 VGND 0.059028f
C3181 a_10108_26262.t2 VGND 0.059028f
C3182 a_10108_26262.n0 VGND 0.136068f
C3183 a_10108_26262.t1 VGND 0.059028f
C3184 a_10108_26262.t0 VGND 0.059028f
C3185 a_10108_26262.n1 VGND 0.258102f
C3186 a_10108_26262.n2 VGND 1.11221f
C3187 a_10108_26262.n3 VGND 0.139449f
C3188 a_10108_26262.t4 VGND 0.059028f
C3189 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3190 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.041341f
C3191 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.096169f
C3192 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3193 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.089265f
C3194 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.083414f
C3195 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3196 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.087824f
C3197 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.03985f
C3198 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3199 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.200787f
C3200 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.202074f
C3201 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C3202 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3203 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3204 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3205 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.107523f
C3206 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3207 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3208 a_10958_37056.t8 VGND 0.024913f
C3209 a_10958_37056.t9 VGND 0.024913f
C3210 a_10958_37056.t6 VGND 0.024913f
C3211 a_10958_37056.n0 VGND 0.059872f
C3212 a_10958_37056.t4 VGND 0.096748f
C3213 a_10958_37056.t2 VGND 0.024913f
C3214 a_10958_37056.t12 VGND 0.024913f
C3215 a_10958_37056.n1 VGND 0.060504f
C3216 a_10958_37056.n2 VGND 0.369187f
C3217 a_10958_37056.t5 VGND 0.024913f
C3218 a_10958_37056.t3 VGND 0.024913f
C3219 a_10958_37056.n3 VGND 0.060504f
C3220 a_10958_37056.n4 VGND 0.182084f
C3221 a_10958_37056.t11 VGND 0.024913f
C3222 a_10958_37056.t1 VGND 0.024913f
C3223 a_10958_37056.n5 VGND 0.060504f
C3224 a_10958_37056.n6 VGND 0.221492f
C3225 a_10958_37056.t7 VGND 0.024913f
C3226 a_10958_37056.t0 VGND 0.024913f
C3227 a_10958_37056.n7 VGND 0.052659f
C3228 a_10958_37056.n8 VGND 0.137512f
C3229 a_10958_37056.n9 VGND 0.342225f
C3230 a_10958_37056.n10 VGND 0.057757f
C3231 a_10958_37056.t10 VGND 0.024913f
C3232 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t7 VGND 0.027086f
C3233 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t3 VGND 0.034765f
C3234 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t5 VGND 0.034765f
C3235 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n0 VGND 0.10415f
C3236 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t0 VGND 0.067642f
C3237 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t1 VGND 0.215011f
C3238 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n1 VGND 0.85898f
C3239 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t4 VGND 0.093153f
C3240 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t2 VGND 0.086397f
C3241 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.t6 VGND 0.093468f
C3242 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n2 VGND 0.091702f
C3243 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n3 VGND 0.063806f
C3244 variable_delay_short_0.variable_delay_unit_5.tristate_inverter_1.en.n4 VGND 0.942937f
C3245 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_1 VGND 0.375772f
C3246 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d VGND 0.696742f
C3247 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 VGND 0.059856f
C3248 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 VGND 0.019094f
C3249 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 VGND 0.041709f
C3250 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 VGND 0.059856f
C3251 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 VGND 0.019094f
C3252 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 VGND 0.04198f
C3253 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 VGND 0.013454f
C3254 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 VGND 0.059856f
C3255 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 VGND 0.019094f
C3256 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 VGND 0.04198f
C3257 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 VGND 0.059856f
C3258 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 VGND 0.019094f
C3259 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 VGND 0.041709f
C3260 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 VGND 0.013307f
C3261 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 VGND 0.351257f
C3262 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 VGND 0.047903f
C3263 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 VGND 0.144997f
C3264 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 VGND 0.368007f
C3265 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 VGND 0.013091f
C3266 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 VGND 0.013091f
C3267 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 VGND 0.030662f
C3268 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 VGND 0.039272f
C3269 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 VGND 0.039272f
C3270 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 VGND 0.080004f
C3271 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 VGND 0.332866f
C3272 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 VGND 0.060722f
C3273 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 VGND 0.060722f
C3274 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 VGND 0.070899f
C3275 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 VGND 0.060722f
C3276 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 VGND 0.060722f
C3277 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 VGND 0.070523f
C3278 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 VGND 0.632153f
C3279 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 VGND 0.045973f
C3280 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 VGND 0.156775f
C3281 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 VGND 0.144997f
C3282 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 VGND 0.240639f
C3283 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 VGND 0.180864f
C3284 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 VGND 0.271416f
C3285 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t3 VGND 0.019446f
C3286 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t6 VGND 0.02496f
C3287 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t2 VGND 0.02496f
C3288 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n0 VGND 0.074774f
C3289 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t1 VGND 0.048564f
C3290 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t0 VGND 0.154367f
C3291 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n1 VGND 0.616703f
C3292 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t7 VGND 0.066879f
C3293 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t5 VGND 0.062029f
C3294 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.t4 VGND 0.067105f
C3295 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n2 VGND 0.065837f
C3296 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n3 VGND 0.045809f
C3297 variable_delay_short_0.variable_delay_unit_3.tristate_inverter_1.en.n4 VGND 0.676981f
C3298 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3299 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.041341f
C3300 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.096169f
C3301 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3302 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.089265f
C3303 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.083414f
C3304 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3305 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.202074f
C3306 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.087824f
C3307 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.03985f
C3308 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3309 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.200787f
C3310 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3311 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.054421f
C3312 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3313 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3314 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.107523f
C3315 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3316 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3317 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3318 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3319 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.087567f
C3320 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.039734f
C3321 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3322 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.089004f
C3323 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.08317f
C3324 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.109331f
C3325 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.041221f
C3326 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.095888f
C3327 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.116125f
C3328 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.108461f
C3329 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.202442f
C3330 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C3331 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.054262f
C3332 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.115417f
C3333 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C3334 a_10108_35390.t0 VGND 0.059028f
C3335 a_10108_35390.t4 VGND 0.059028f
C3336 a_10108_35390.t3 VGND 0.059028f
C3337 a_10108_35390.n0 VGND 0.136068f
C3338 a_10108_35390.t2 VGND 0.059028f
C3339 a_10108_35390.t5 VGND 0.059028f
C3340 a_10108_35390.n1 VGND 0.258102f
C3341 a_10108_35390.n2 VGND 1.11221f
C3342 a_10108_35390.n3 VGND 0.139449f
C3343 a_10108_35390.t1 VGND 0.059028f
C3344 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3345 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3346 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.087567f
C3347 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.039734f
C3348 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3349 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C3350 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C3351 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.054262f
C3352 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.115417f
C3353 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.089004f
C3354 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.08317f
C3355 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C3356 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.041221f
C3357 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.095888f
C3358 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C3359 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.108461f
C3360 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C3361 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3362 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.041341f
C3363 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.096169f
C3364 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3365 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.089265f
C3366 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.083414f
C3367 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3368 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.202074f
C3369 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.087824f
C3370 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C3371 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3372 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.200787f
C3373 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.054421f
C3374 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3375 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3376 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3377 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.107523f
C3378 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3379 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3380 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3381 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3382 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.087567f
C3383 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.039734f
C3384 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3385 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.202442f
C3386 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.054262f
C3387 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C3388 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.115417f
C3389 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.089004f
C3390 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.08317f
C3391 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.109331f
C3392 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.041221f
C3393 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.095888f
C3394 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.116125f
C3395 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.108461f
C3396 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.202442f
C3397 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t3 VGND 0.019446f
C3398 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t5 VGND 0.02496f
C3399 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t7 VGND 0.02496f
C3400 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n0 VGND 0.074774f
C3401 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t1 VGND 0.048564f
C3402 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t0 VGND 0.154367f
C3403 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n1 VGND 0.616703f
C3404 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t6 VGND 0.066879f
C3405 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t4 VGND 0.062029f
C3406 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.t2 VGND 0.067105f
C3407 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n2 VGND 0.065837f
C3408 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n3 VGND 0.045809f
C3409 variable_delay_short_0.variable_delay_unit_0.tristate_inverter_1.en.n4 VGND 0.676981f
C3410 a_10958_23364.t5 VGND 0.024913f
C3411 a_10958_23364.t1 VGND 0.096748f
C3412 a_10958_23364.t10 VGND 0.024913f
C3413 a_10958_23364.t11 VGND 0.024913f
C3414 a_10958_23364.n0 VGND 0.060504f
C3415 a_10958_23364.n1 VGND 0.369187f
C3416 a_10958_23364.t12 VGND 0.024913f
C3417 a_10958_23364.t9 VGND 0.024913f
C3418 a_10958_23364.n2 VGND 0.060504f
C3419 a_10958_23364.n3 VGND 0.182084f
C3420 a_10958_23364.t8 VGND 0.024913f
C3421 a_10958_23364.t0 VGND 0.024913f
C3422 a_10958_23364.n4 VGND 0.060504f
C3423 a_10958_23364.n5 VGND 0.221492f
C3424 a_10958_23364.t2 VGND 0.024913f
C3425 a_10958_23364.t7 VGND 0.024913f
C3426 a_10958_23364.n6 VGND 0.052659f
C3427 a_10958_23364.n7 VGND 0.137512f
C3428 a_10958_23364.t3 VGND 0.024913f
C3429 a_10958_23364.t4 VGND 0.024913f
C3430 a_10958_23364.n8 VGND 0.057757f
C3431 a_10958_23364.n9 VGND 0.342225f
C3432 a_10958_23364.n10 VGND 0.059872f
C3433 a_10958_23364.t6 VGND 0.024913f
C3434 a_10108_28544.t0 VGND 0.059028f
C3435 a_10108_28544.t3 VGND 0.059028f
C3436 a_10108_28544.t5 VGND 0.059028f
C3437 a_10108_28544.n0 VGND 0.136068f
C3438 a_10108_28544.t4 VGND 0.059028f
C3439 a_10108_28544.t2 VGND 0.059028f
C3440 a_10108_28544.n1 VGND 0.258102f
C3441 a_10108_28544.n2 VGND 1.11221f
C3442 a_10108_28544.n3 VGND 0.139449f
C3443 a_10108_28544.t1 VGND 0.059028f
C3444 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 VGND 1.51406f
C3445 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 VGND 0.930597f
C3446 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 VGND 0.087567f
C3447 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 VGND 0.039734f
C3448 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 VGND 0.097942f
C3449 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 VGND 0.202442f
C3450 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 VGND 0.089004f
C3451 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 VGND 0.08317f
C3452 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 VGND 0.109331f
C3453 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 VGND 0.041221f
C3454 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 VGND 0.095888f
C3455 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 VGND 0.116125f
C3456 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 VGND 0.108461f
C3457 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 VGND 0.202442f
C3458 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 VGND 0.054262f
C3459 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 VGND 0.054262f
C3460 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 VGND 0.115417f
C3461 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3462 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.041341f
C3463 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.096169f
C3464 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3465 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.089265f
C3466 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.083414f
C3467 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3468 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.087824f
C3469 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C3470 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3471 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.200787f
C3472 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.202074f
C3473 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.054421f
C3474 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.054421f
C3475 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3476 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3477 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.107523f
C3478 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3479 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3480 a_10958_39338.t3 VGND 0.024913f
C3481 a_10958_39338.t1 VGND 0.096748f
C3482 a_10958_39338.t8 VGND 0.024913f
C3483 a_10958_39338.t0 VGND 0.024913f
C3484 a_10958_39338.n0 VGND 0.060504f
C3485 a_10958_39338.n1 VGND 0.369187f
C3486 a_10958_39338.t12 VGND 0.024913f
C3487 a_10958_39338.t11 VGND 0.024913f
C3488 a_10958_39338.n2 VGND 0.060504f
C3489 a_10958_39338.n3 VGND 0.182084f
C3490 a_10958_39338.t9 VGND 0.024913f
C3491 a_10958_39338.t7 VGND 0.024913f
C3492 a_10958_39338.n4 VGND 0.060504f
C3493 a_10958_39338.n5 VGND 0.221492f
C3494 a_10958_39338.t2 VGND 0.024913f
C3495 a_10958_39338.t10 VGND 0.024913f
C3496 a_10958_39338.n6 VGND 0.052659f
C3497 a_10958_39338.n7 VGND 0.137512f
C3498 a_10958_39338.t4 VGND 0.024913f
C3499 a_10958_39338.t5 VGND 0.024913f
C3500 a_10958_39338.n8 VGND 0.057757f
C3501 a_10958_39338.n9 VGND 0.342225f
C3502 a_10958_39338.n10 VGND 0.059872f
C3503 a_10958_39338.t6 VGND 0.024913f
C3504 a_10108_39954.t1 VGND 0.059028f
C3505 a_10108_39954.t3 VGND 0.059028f
C3506 a_10108_39954.t2 VGND 0.059028f
C3507 a_10108_39954.n0 VGND 0.136068f
C3508 a_10108_39954.t4 VGND 0.059028f
C3509 a_10108_39954.t5 VGND 0.059028f
C3510 a_10108_39954.n1 VGND 0.258102f
C3511 a_10108_39954.n2 VGND 1.11221f
C3512 a_10108_39954.n3 VGND 0.139449f
C3513 a_10108_39954.t0 VGND 0.059028f
C3514 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd VGND 0.503525f
C3515 tdc_0.vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 VGND 0.130197f
C3516 tdc_0.vernier_delay_line_0.delay_unit_2_0.in_2 VGND 0.189073f
C3517 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 VGND 0.09757f
C3518 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 VGND 0.030153f
C3519 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 VGND 0.265657f
C3520 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 VGND 0.039259f
C3521 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 VGND 0.012524f
C3522 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 VGND 0.027534f
C3523 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 VGND 0.039259f
C3524 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 VGND 0.012524f
C3525 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 VGND 0.027357f
C3526 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 VGND 0.008823f
C3527 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 VGND 0.039259f
C3528 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 VGND 0.012524f
C3529 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 VGND 0.027534f
C3530 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 VGND 0.039259f
C3531 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 VGND 0.012524f
C3532 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 VGND 0.027357f
C3533 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 VGND 0.008728f
C3534 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 VGND 0.135162f
C3535 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 VGND 0.046129f
C3536 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 VGND 0.046129f
C3537 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 VGND 0.054044f
C3538 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 VGND 0.046129f
C3539 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 VGND 0.046129f
C3540 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 VGND 0.0538f
C3541 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 VGND 0.495704f
C3542 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 VGND 0.025758f
C3543 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 VGND 0.025758f
C3544 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 VGND 0.055083f
C3545 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 VGND 0.008586f
C3546 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 VGND 0.008586f
C3547 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 VGND 0.01864f
C3548 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 VGND 0.221512f
C3549 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 VGND 0.09757f
C3550 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 VGND 0.030153f
C3551 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 VGND 0.234486f
C3552 tdc_0.vernier_delay_line_0.stop_strong.t78 VGND 0.078403f
C3553 tdc_0.vernier_delay_line_0.stop_strong.t43 VGND 0.073263f
C3554 tdc_0.vernier_delay_line_0.stop_strong.n0 VGND 0.070349f
C3555 tdc_0.vernier_delay_line_0.stop_strong.t55 VGND 0.073263f
C3556 tdc_0.vernier_delay_line_0.stop_strong.n1 VGND 0.040134f
C3557 tdc_0.vernier_delay_line_0.stop_strong.t72 VGND 0.073263f
C3558 tdc_0.vernier_delay_line_0.stop_strong.n2 VGND 0.040134f
C3559 tdc_0.vernier_delay_line_0.stop_strong.t37 VGND 0.073263f
C3560 tdc_0.vernier_delay_line_0.stop_strong.n3 VGND 0.064514f
C3561 tdc_0.vernier_delay_line_0.stop_strong.t56 VGND 0.093756f
C3562 tdc_0.vernier_delay_line_0.stop_strong.t87 VGND 0.093545f
C3563 tdc_0.vernier_delay_line_0.stop_strong.n4 VGND 0.403473f
C3564 tdc_0.vernier_delay_line_0.stop_strong.n5 VGND 0.933667f
C3565 tdc_0.vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk VGND 1.3151f
C3566 tdc_0.vernier_delay_line_0.stop_strong.t67 VGND 0.078403f
C3567 tdc_0.vernier_delay_line_0.stop_strong.t33 VGND 0.073263f
C3568 tdc_0.vernier_delay_line_0.stop_strong.n6 VGND 0.070349f
C3569 tdc_0.vernier_delay_line_0.stop_strong.t60 VGND 0.073263f
C3570 tdc_0.vernier_delay_line_0.stop_strong.n7 VGND 0.040134f
C3571 tdc_0.vernier_delay_line_0.stop_strong.t82 VGND 0.073263f
C3572 tdc_0.vernier_delay_line_0.stop_strong.n8 VGND 0.040134f
C3573 tdc_0.vernier_delay_line_0.stop_strong.t46 VGND 0.073263f
C3574 tdc_0.vernier_delay_line_0.stop_strong.n9 VGND 0.064514f
C3575 tdc_0.vernier_delay_line_0.stop_strong.t80 VGND 0.093756f
C3576 tdc_0.vernier_delay_line_0.stop_strong.t39 VGND 0.093545f
C3577 tdc_0.vernier_delay_line_0.stop_strong.n10 VGND 0.403473f
C3578 tdc_0.vernier_delay_line_0.stop_strong.n11 VGND 0.777822f
C3579 tdc_0.vernier_delay_line_0.stop_strong.n12 VGND 0.697925f
C3580 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3581 tdc_0.vernier_delay_line_0.stop_strong.t52 VGND 0.078403f
C3582 tdc_0.vernier_delay_line_0.stop_strong.t68 VGND 0.073263f
C3583 tdc_0.vernier_delay_line_0.stop_strong.n13 VGND 0.070349f
C3584 tdc_0.vernier_delay_line_0.stop_strong.t35 VGND 0.073263f
C3585 tdc_0.vernier_delay_line_0.stop_strong.n14 VGND 0.040134f
C3586 tdc_0.vernier_delay_line_0.stop_strong.t51 VGND 0.073263f
C3587 tdc_0.vernier_delay_line_0.stop_strong.n15 VGND 0.040134f
C3588 tdc_0.vernier_delay_line_0.stop_strong.t64 VGND 0.073263f
C3589 tdc_0.vernier_delay_line_0.stop_strong.n16 VGND 0.064514f
C3590 tdc_0.vernier_delay_line_0.stop_strong.t61 VGND 0.093756f
C3591 tdc_0.vernier_delay_line_0.stop_strong.t59 VGND 0.093545f
C3592 tdc_0.vernier_delay_line_0.stop_strong.n17 VGND 0.403473f
C3593 tdc_0.vernier_delay_line_0.stop_strong.n18 VGND 0.777822f
C3594 tdc_0.vernier_delay_line_0.stop_strong.n19 VGND 0.697925f
C3595 tdc_0.vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3596 tdc_0.vernier_delay_line_0.stop_strong.t40 VGND 0.078403f
C3597 tdc_0.vernier_delay_line_0.stop_strong.t53 VGND 0.073263f
C3598 tdc_0.vernier_delay_line_0.stop_strong.n20 VGND 0.070349f
C3599 tdc_0.vernier_delay_line_0.stop_strong.t69 VGND 0.073263f
C3600 tdc_0.vernier_delay_line_0.stop_strong.n21 VGND 0.040134f
C3601 tdc_0.vernier_delay_line_0.stop_strong.t71 VGND 0.073263f
C3602 tdc_0.vernier_delay_line_0.stop_strong.n22 VGND 0.040134f
C3603 tdc_0.vernier_delay_line_0.stop_strong.t36 VGND 0.073263f
C3604 tdc_0.vernier_delay_line_0.stop_strong.n23 VGND 0.064514f
C3605 tdc_0.vernier_delay_line_0.stop_strong.t49 VGND 0.093756f
C3606 tdc_0.vernier_delay_line_0.stop_strong.t45 VGND 0.093545f
C3607 tdc_0.vernier_delay_line_0.stop_strong.n24 VGND 0.403473f
C3608 tdc_0.vernier_delay_line_0.stop_strong.n25 VGND 0.777822f
C3609 tdc_0.vernier_delay_line_0.stop_strong.n26 VGND 0.697925f
C3610 tdc_0.vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3611 tdc_0.vernier_delay_line_0.stop_strong.t70 VGND 0.078403f
C3612 tdc_0.vernier_delay_line_0.stop_strong.t42 VGND 0.073263f
C3613 tdc_0.vernier_delay_line_0.stop_strong.n27 VGND 0.070349f
C3614 tdc_0.vernier_delay_line_0.stop_strong.t44 VGND 0.073263f
C3615 tdc_0.vernier_delay_line_0.stop_strong.n28 VGND 0.040134f
C3616 tdc_0.vernier_delay_line_0.stop_strong.t57 VGND 0.073263f
C3617 tdc_0.vernier_delay_line_0.stop_strong.n29 VGND 0.040134f
C3618 tdc_0.vernier_delay_line_0.stop_strong.t73 VGND 0.073263f
C3619 tdc_0.vernier_delay_line_0.stop_strong.n30 VGND 0.064514f
C3620 tdc_0.vernier_delay_line_0.stop_strong.t66 VGND 0.093756f
C3621 tdc_0.vernier_delay_line_0.stop_strong.t77 VGND 0.093545f
C3622 tdc_0.vernier_delay_line_0.stop_strong.n31 VGND 0.403473f
C3623 tdc_0.vernier_delay_line_0.stop_strong.n32 VGND 0.777822f
C3624 tdc_0.vernier_delay_line_0.stop_strong.n33 VGND 0.697925f
C3625 tdc_0.vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3626 tdc_0.vernier_delay_line_0.stop_strong.t81 VGND 0.078403f
C3627 tdc_0.vernier_delay_line_0.stop_strong.t83 VGND 0.073263f
C3628 tdc_0.vernier_delay_line_0.stop_strong.n34 VGND 0.070349f
C3629 tdc_0.vernier_delay_line_0.stop_strong.t47 VGND 0.073263f
C3630 tdc_0.vernier_delay_line_0.stop_strong.n35 VGND 0.040134f
C3631 tdc_0.vernier_delay_line_0.stop_strong.t62 VGND 0.073263f
C3632 tdc_0.vernier_delay_line_0.stop_strong.n36 VGND 0.040134f
C3633 tdc_0.vernier_delay_line_0.stop_strong.t84 VGND 0.073263f
C3634 tdc_0.vernier_delay_line_0.stop_strong.n37 VGND 0.064514f
C3635 tdc_0.vernier_delay_line_0.stop_strong.t76 VGND 0.093756f
C3636 tdc_0.vernier_delay_line_0.stop_strong.t74 VGND 0.093545f
C3637 tdc_0.vernier_delay_line_0.stop_strong.n38 VGND 0.403473f
C3638 tdc_0.vernier_delay_line_0.stop_strong.n39 VGND 0.777822f
C3639 tdc_0.vernier_delay_line_0.stop_strong.n40 VGND 0.697925f
C3640 tdc_0.vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3641 tdc_0.vernier_delay_line_0.stop_strong.t38 VGND 0.078403f
C3642 tdc_0.vernier_delay_line_0.stop_strong.t65 VGND 0.073263f
C3643 tdc_0.vernier_delay_line_0.stop_strong.n41 VGND 0.070349f
C3644 tdc_0.vernier_delay_line_0.stop_strong.t85 VGND 0.073263f
C3645 tdc_0.vernier_delay_line_0.stop_strong.n42 VGND 0.040134f
C3646 tdc_0.vernier_delay_line_0.stop_strong.t50 VGND 0.073263f
C3647 tdc_0.vernier_delay_line_0.stop_strong.n43 VGND 0.040134f
C3648 tdc_0.vernier_delay_line_0.stop_strong.t63 VGND 0.073263f
C3649 tdc_0.vernier_delay_line_0.stop_strong.n44 VGND 0.064514f
C3650 tdc_0.vernier_delay_line_0.stop_strong.t48 VGND 0.093756f
C3651 tdc_0.vernier_delay_line_0.stop_strong.t58 VGND 0.093545f
C3652 tdc_0.vernier_delay_line_0.stop_strong.n45 VGND 0.403473f
C3653 tdc_0.vernier_delay_line_0.stop_strong.n46 VGND 0.777822f
C3654 tdc_0.vernier_delay_line_0.stop_strong.n47 VGND 0.697925f
C3655 tdc_0.vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk VGND 0.626873f
C3656 tdc_0.vernier_delay_line_0.stop_strong.t75 VGND 0.078403f
C3657 tdc_0.vernier_delay_line_0.stop_strong.t41 VGND 0.073263f
C3658 tdc_0.vernier_delay_line_0.stop_strong.n48 VGND 0.070349f
C3659 tdc_0.vernier_delay_line_0.stop_strong.t54 VGND 0.073263f
C3660 tdc_0.vernier_delay_line_0.stop_strong.n49 VGND 0.040134f
C3661 tdc_0.vernier_delay_line_0.stop_strong.t32 VGND 0.073263f
C3662 tdc_0.vernier_delay_line_0.stop_strong.n50 VGND 0.040134f
C3663 tdc_0.vernier_delay_line_0.stop_strong.t34 VGND 0.073263f
C3664 tdc_0.vernier_delay_line_0.stop_strong.n51 VGND 0.064514f
C3665 tdc_0.vernier_delay_line_0.stop_strong.t86 VGND 0.093756f
C3666 tdc_0.vernier_delay_line_0.stop_strong.t79 VGND 0.093545f
C3667 tdc_0.vernier_delay_line_0.stop_strong.n52 VGND 0.403473f
C3668 tdc_0.vernier_delay_line_0.stop_strong.n53 VGND 0.777822f
C3669 tdc_0.vernier_delay_line_0.stop_strong.n54 VGND 0.697925f
C3670 tdc_0.vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk VGND 0.971005f
C3671 tdc_0.vernier_delay_line_0.stop_strong.t27 VGND 0.181057f
C3672 tdc_0.vernier_delay_line_0.stop_strong.t13 VGND 0.055955f
C3673 tdc_0.vernier_delay_line_0.stop_strong.n55 VGND 0.420822f
C3674 tdc_0.vernier_delay_line_0.stop_strong.t20 VGND 0.181057f
C3675 tdc_0.vernier_delay_line_0.stop_strong.t6 VGND 0.055955f
C3676 tdc_0.vernier_delay_line_0.stop_strong.n56 VGND 0.413796f
C3677 tdc_0.vernier_delay_line_0.stop_strong.n57 VGND 0.17535f
C3678 tdc_0.vernier_delay_line_0.stop_strong.t30 VGND 0.181057f
C3679 tdc_0.vernier_delay_line_0.stop_strong.t0 VGND 0.055955f
C3680 tdc_0.vernier_delay_line_0.stop_strong.n58 VGND 0.413796f
C3681 tdc_0.vernier_delay_line_0.stop_strong.n59 VGND 0.11234f
C3682 tdc_0.vernier_delay_line_0.stop_strong.t23 VGND 0.181057f
C3683 tdc_0.vernier_delay_line_0.stop_strong.t9 VGND 0.055955f
C3684 tdc_0.vernier_delay_line_0.stop_strong.n60 VGND 0.413796f
C3685 tdc_0.vernier_delay_line_0.stop_strong.n61 VGND 0.11234f
C3686 tdc_0.vernier_delay_line_0.stop_strong.t17 VGND 0.181057f
C3687 tdc_0.vernier_delay_line_0.stop_strong.t3 VGND 0.055955f
C3688 tdc_0.vernier_delay_line_0.stop_strong.n62 VGND 0.413796f
C3689 tdc_0.vernier_delay_line_0.stop_strong.n63 VGND 0.11234f
C3690 tdc_0.vernier_delay_line_0.stop_strong.t26 VGND 0.181057f
C3691 tdc_0.vernier_delay_line_0.stop_strong.t12 VGND 0.055955f
C3692 tdc_0.vernier_delay_line_0.stop_strong.n64 VGND 0.413796f
C3693 tdc_0.vernier_delay_line_0.stop_strong.n65 VGND 0.11234f
C3694 tdc_0.vernier_delay_line_0.stop_strong.t16 VGND 0.181057f
C3695 tdc_0.vernier_delay_line_0.stop_strong.t2 VGND 0.055955f
C3696 tdc_0.vernier_delay_line_0.stop_strong.n66 VGND 0.413796f
C3697 tdc_0.vernier_delay_line_0.stop_strong.n67 VGND 0.11234f
C3698 tdc_0.vernier_delay_line_0.stop_strong.t25 VGND 0.181057f
C3699 tdc_0.vernier_delay_line_0.stop_strong.t11 VGND 0.055955f
C3700 tdc_0.vernier_delay_line_0.stop_strong.n68 VGND 0.413796f
C3701 tdc_0.vernier_delay_line_0.stop_strong.n69 VGND 0.11234f
C3702 tdc_0.vernier_delay_line_0.stop_strong.t19 VGND 0.181057f
C3703 tdc_0.vernier_delay_line_0.stop_strong.t5 VGND 0.055955f
C3704 tdc_0.vernier_delay_line_0.stop_strong.n70 VGND 0.413796f
C3705 tdc_0.vernier_delay_line_0.stop_strong.n71 VGND 0.11234f
C3706 tdc_0.vernier_delay_line_0.stop_strong.t29 VGND 0.181057f
C3707 tdc_0.vernier_delay_line_0.stop_strong.t15 VGND 0.055955f
C3708 tdc_0.vernier_delay_line_0.stop_strong.n72 VGND 0.413796f
C3709 tdc_0.vernier_delay_line_0.stop_strong.n73 VGND 0.11234f
C3710 tdc_0.vernier_delay_line_0.stop_strong.t22 VGND 0.181057f
C3711 tdc_0.vernier_delay_line_0.stop_strong.t8 VGND 0.055955f
C3712 tdc_0.vernier_delay_line_0.stop_strong.n74 VGND 0.413796f
C3713 tdc_0.vernier_delay_line_0.stop_strong.n75 VGND 0.11234f
C3714 tdc_0.vernier_delay_line_0.stop_strong.t24 VGND 0.181057f
C3715 tdc_0.vernier_delay_line_0.stop_strong.t10 VGND 0.055955f
C3716 tdc_0.vernier_delay_line_0.stop_strong.n76 VGND 0.413796f
C3717 tdc_0.vernier_delay_line_0.stop_strong.n77 VGND 0.11234f
C3718 tdc_0.vernier_delay_line_0.stop_strong.t18 VGND 0.181057f
C3719 tdc_0.vernier_delay_line_0.stop_strong.t4 VGND 0.055955f
C3720 tdc_0.vernier_delay_line_0.stop_strong.n78 VGND 0.413796f
C3721 tdc_0.vernier_delay_line_0.stop_strong.n79 VGND 0.11234f
C3722 tdc_0.vernier_delay_line_0.stop_strong.t28 VGND 0.181057f
C3723 tdc_0.vernier_delay_line_0.stop_strong.t14 VGND 0.055955f
C3724 tdc_0.vernier_delay_line_0.stop_strong.n80 VGND 0.413796f
C3725 tdc_0.vernier_delay_line_0.stop_strong.n81 VGND 0.11234f
C3726 tdc_0.vernier_delay_line_0.stop_strong.t21 VGND 0.181057f
C3727 tdc_0.vernier_delay_line_0.stop_strong.t7 VGND 0.055955f
C3728 tdc_0.vernier_delay_line_0.stop_strong.n82 VGND 0.413796f
C3729 tdc_0.vernier_delay_line_0.stop_strong.n83 VGND 0.110532f
C3730 tdc_0.vernier_delay_line_0.stop_strong.n84 VGND 1.2768f
C3731 tdc_0.vernier_delay_line_0.stop_strong.t1 VGND 0.055955f
C3732 tdc_0.vernier_delay_line_0.stop_strong.n85 VGND 0.097761f
C3733 tdc_0.vernier_delay_line_0.stop_strong.t31 VGND 0.179153f
C3734 tdc_0.vernier_delay_line_0.stop_strong.n86 VGND 0.326098f
C3735 tdc_0.stop_buffer_0.stop_strong VGND 0.031003f
C3736 a_9330_16954.t4 VGND 0.228995f
C3737 a_9330_16954.t17 VGND 0.093349f
C3738 a_9330_16954.t13 VGND 0.030133f
C3739 a_9330_16954.n0 VGND 0.086421f
C3740 a_9330_16954.t9 VGND 0.093349f
C3741 a_9330_16954.t38 VGND 0.030133f
C3742 a_9330_16954.n1 VGND 0.088816f
C3743 a_9330_16954.t29 VGND 0.093349f
C3744 a_9330_16954.t26 VGND 0.030133f
C3745 a_9330_16954.n2 VGND 0.088354f
C3746 a_9330_16954.n3 VGND 0.389976f
C3747 a_9330_16954.t16 VGND 0.093349f
C3748 a_9330_16954.t12 VGND 0.030133f
C3749 a_9330_16954.n4 VGND 0.088354f
C3750 a_9330_16954.n5 VGND 0.217864f
C3751 a_9330_16954.t35 VGND 0.093349f
C3752 a_9330_16954.t32 VGND 0.030133f
C3753 a_9330_16954.n6 VGND 0.088354f
C3754 a_9330_16954.n7 VGND 0.217864f
C3755 a_9330_16954.t23 VGND 0.093349f
C3756 a_9330_16954.t20 VGND 0.030133f
C3757 a_9330_16954.n8 VGND 0.088354f
C3758 a_9330_16954.n9 VGND 0.217864f
C3759 a_9330_16954.t25 VGND 0.093349f
C3760 a_9330_16954.t22 VGND 0.030133f
C3761 a_9330_16954.n10 VGND 0.088354f
C3762 a_9330_16954.n11 VGND 0.217864f
C3763 a_9330_16954.t11 VGND 0.093349f
C3764 a_9330_16954.t8 VGND 0.030133f
C3765 a_9330_16954.n12 VGND 0.088354f
C3766 a_9330_16954.n13 VGND 0.217864f
C3767 a_9330_16954.t31 VGND 0.093349f
C3768 a_9330_16954.t28 VGND 0.030133f
C3769 a_9330_16954.n14 VGND 0.088354f
C3770 a_9330_16954.n15 VGND 0.217864f
C3771 a_9330_16954.t19 VGND 0.093349f
C3772 a_9330_16954.t15 VGND 0.030133f
C3773 a_9330_16954.n16 VGND 0.088354f
C3774 a_9330_16954.n17 VGND 0.217864f
C3775 a_9330_16954.t37 VGND 0.093349f
C3776 a_9330_16954.t34 VGND 0.030133f
C3777 a_9330_16954.n18 VGND 0.088354f
C3778 a_9330_16954.n19 VGND 0.217864f
C3779 a_9330_16954.t18 VGND 0.093349f
C3780 a_9330_16954.t14 VGND 0.030133f
C3781 a_9330_16954.n20 VGND 0.088354f
C3782 a_9330_16954.n21 VGND 0.217864f
C3783 a_9330_16954.t36 VGND 0.093349f
C3784 a_9330_16954.t33 VGND 0.030133f
C3785 a_9330_16954.n22 VGND 0.088354f
C3786 a_9330_16954.n23 VGND 0.217864f
C3787 a_9330_16954.t24 VGND 0.093349f
C3788 a_9330_16954.t21 VGND 0.030133f
C3789 a_9330_16954.n24 VGND 0.088354f
C3790 a_9330_16954.n25 VGND 0.217864f
C3791 a_9330_16954.t10 VGND 0.093349f
C3792 a_9330_16954.t39 VGND 0.030133f
C3793 a_9330_16954.n26 VGND 0.088354f
C3794 a_9330_16954.n27 VGND 0.217864f
C3795 a_9330_16954.t30 VGND 0.093349f
C3796 a_9330_16954.t27 VGND 0.030133f
C3797 a_9330_16954.n28 VGND 0.088354f
C3798 a_9330_16954.n29 VGND 0.289551f
C3799 a_9330_16954.n30 VGND 0.109352f
C3800 a_9330_16954.n31 VGND 0.42154f
C3801 a_9330_16954.t0 VGND 0.071536f
C3802 a_9330_16954.n32 VGND 0.133321f
C3803 a_9330_16954.t6 VGND 0.231476f
C3804 a_9330_16954.t2 VGND 0.071536f
C3805 a_9330_16954.n33 VGND 0.529025f
C3806 a_9330_16954.n34 VGND 0.22418f
C3807 a_9330_16954.t5 VGND 0.231476f
C3808 a_9330_16954.t1 VGND 0.071536f
C3809 a_9330_16954.n35 VGND 0.538008f
C3810 a_9330_16954.n36 VGND 0.22418f
C3811 a_9330_16954.t3 VGND 0.071536f
C3812 a_9330_16954.n37 VGND 0.529025f
C3813 a_9330_16954.t7 VGND 0.231476f
C3814 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 VGND 1.05156f
C3815 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 VGND 0.041341f
C3816 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 VGND 0.096169f
C3817 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 VGND 0.116334f
C3818 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 VGND 0.089265f
C3819 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 VGND 0.083414f
C3820 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 VGND 0.110889f
C3821 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 VGND 0.202074f
C3822 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 VGND 0.087824f
C3823 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 VGND 0.03985f
C3824 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 VGND 0.098113f
C3825 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 VGND 0.200787f
C3826 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 VGND 0.054421f
C3827 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 VGND 0.054421f
C3828 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 VGND 0.114315f
C3829 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 VGND 0.385552f
C3830 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 VGND 0.107523f
C3831 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 VGND 0.139754f
C3832 tdc_0.vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 VGND 1.24397f
C3833 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t3 VGND 0.019446f
C3834 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t5 VGND 0.02496f
C3835 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t7 VGND 0.02496f
C3836 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n0 VGND 0.074774f
C3837 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t1 VGND 0.048564f
C3838 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t0 VGND 0.154367f
C3839 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n1 VGND 0.616703f
C3840 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t6 VGND 0.066879f
C3841 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t4 VGND 0.062029f
C3842 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.t2 VGND 0.067105f
C3843 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n2 VGND 0.065837f
C3844 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n3 VGND 0.045809f
C3845 variable_delay_short_0.variable_delay_unit_1.tristate_inverter_1.en.n4 VGND 0.676981f
C3846 tdc_0.start_buffer_0.start_delay.t8 VGND 0.069408f
C3847 tdc_0.start_buffer_0.start_delay.t15 VGND 0.022142f
C3848 tdc_0.start_buffer_0.start_delay.n0 VGND 0.04868f
C3849 tdc_0.start_buffer_0.start_delay.t14 VGND 0.069408f
C3850 tdc_0.start_buffer_0.start_delay.t12 VGND 0.022142f
C3851 tdc_0.start_buffer_0.start_delay.n1 VGND 0.048366f
C3852 tdc_0.start_buffer_0.start_delay.n2 VGND 0.015598f
C3853 tdc_0.start_buffer_0.start_delay.t13 VGND 0.069408f
C3854 tdc_0.start_buffer_0.start_delay.t11 VGND 0.022142f
C3855 tdc_0.start_buffer_0.start_delay.n3 VGND 0.04868f
C3856 tdc_0.start_buffer_0.start_delay.t10 VGND 0.069408f
C3857 tdc_0.start_buffer_0.start_delay.t9 VGND 0.022142f
C3858 tdc_0.start_buffer_0.start_delay.n4 VGND 0.048366f
C3859 tdc_0.start_buffer_0.start_delay.n5 VGND 0.015431f
C3860 tdc_0.start_buffer_0.start_delay.n6 VGND 0.181697f
C3861 tdc_0.start_buffer_0.start_delay.t5 VGND 0.1725f
C3862 tdc_0.start_buffer_0.start_delay.t0 VGND 0.05331f
C3863 tdc_0.start_buffer_0.start_delay.n7 VGND 0.471528f
C3864 tdc_0.start_buffer_0.start_delay.t6 VGND 0.1725f
C3865 tdc_0.start_buffer_0.start_delay.t1 VGND 0.05331f
C3866 tdc_0.start_buffer_0.start_delay.n8 VGND 0.400932f
C3867 tdc_0.start_buffer_0.start_delay.t4 VGND 0.1725f
C3868 tdc_0.start_buffer_0.start_delay.t7 VGND 0.05331f
C3869 tdc_0.start_buffer_0.start_delay.n9 VGND 0.394238f
C3870 tdc_0.start_buffer_0.start_delay.n10 VGND 0.167063f
C3871 tdc_0.start_buffer_0.start_delay.t3 VGND 0.170686f
C3872 tdc_0.start_buffer_0.start_delay.n11 VGND 0.310685f
C3873 tdc_0.start_buffer_0.start_delay.t2 VGND 0.05331f
C3874 tdc_0.start_buffer_0.start_delay.n12 VGND 0.09314f
C3875 tdc_0.start_buffer_0.start_delay.n13 VGND 0.131763f
C3876 tdc_0.start_buffer_0.start_delay.n14 VGND 0.129117f
C3877 tdc_0.start_buffer_0.start_buff.t15 VGND 0.079205f
C3878 tdc_0.start_buffer_0.start_buff.t12 VGND 0.025267f
C3879 tdc_0.start_buffer_0.start_buff.n0 VGND 0.055193f
C3880 tdc_0.start_buffer_0.start_buff.t11 VGND 0.079205f
C3881 tdc_0.start_buffer_0.start_buff.t20 VGND 0.025267f
C3882 tdc_0.start_buffer_0.start_buff.n1 VGND 0.055551f
C3883 tdc_0.start_buffer_0.start_buff.n2 VGND 0.017803f
C3884 tdc_0.start_buffer_0.start_buff.t19 VGND 0.079205f
C3885 tdc_0.start_buffer_0.start_buff.t17 VGND 0.025267f
C3886 tdc_0.start_buffer_0.start_buff.n3 VGND 0.055551f
C3887 tdc_0.start_buffer_0.start_buff.t13 VGND 0.079205f
C3888 tdc_0.start_buffer_0.start_buff.t23 VGND 0.025267f
C3889 tdc_0.start_buffer_0.start_buff.n4 VGND 0.055193f
C3890 tdc_0.start_buffer_0.start_buff.n5 VGND 0.017609f
C3891 tdc_0.start_buffer_0.start_buff.n6 VGND 0.464807f
C3892 tdc_0.start_buffer_0.start_buff.t9 VGND 0.063388f
C3893 tdc_0.start_buffer_0.start_buff.t8 VGND 0.19187f
C3894 tdc_0.start_buffer_0.start_buff.n7 VGND 0.486972f
C3895 tdc_0.start_buffer_0.start_buff.n8 VGND 0.25373f
C3896 tdc_0.start_buffer_0.start_buff.t5 VGND 0.19187f
C3897 tdc_0.start_buffer_0.start_buff.n9 VGND 0.435589f
C3898 tdc_0.start_buffer_0.start_buff.t10 VGND 0.079384f
C3899 tdc_0.start_buffer_0.start_buff.t22 VGND 0.025625f
C3900 tdc_0.start_buffer_0.start_buff.n10 VGND 0.073493f
C3901 tdc_0.start_buffer_0.start_buff.t21 VGND 0.079384f
C3902 tdc_0.start_buffer_0.start_buff.t18 VGND 0.025625f
C3903 tdc_0.start_buffer_0.start_buff.n11 VGND 0.07553f
C3904 tdc_0.start_buffer_0.start_buff.t16 VGND 0.079384f
C3905 tdc_0.start_buffer_0.start_buff.t14 VGND 0.025625f
C3906 tdc_0.start_buffer_0.start_buff.n12 VGND 0.075137f
C3907 tdc_0.start_buffer_0.start_buff.n13 VGND 0.3926f
C3908 tdc_0.start_buffer_0.start_buff.n14 VGND 0.092517f
C3909 tdc_0.start_buffer_0.start_buff.n15 VGND 0.090637f
C3910 tdc_0.start_buffer_0.start_buff.t1 VGND 0.060835f
C3911 tdc_0.start_buffer_0.start_buff.n16 VGND 0.10659f
C3912 tdc_0.start_buffer_0.start_buff.t6 VGND 0.196849f
C3913 tdc_0.start_buffer_0.start_buff.t2 VGND 0.060835f
C3914 tdc_0.start_buffer_0.start_buff.n17 VGND 0.457525f
C3915 tdc_0.start_buffer_0.start_buff.t4 VGND 0.196849f
C3916 tdc_0.start_buffer_0.start_buff.t0 VGND 0.060835f
C3917 tdc_0.start_buffer_0.start_buff.n18 VGND 0.449886f
C3918 tdc_0.start_buffer_0.start_buff.n19 VGND 0.190644f
C3919 tdc_0.start_buffer_0.start_buff.t7 VGND 0.196849f
C3920 tdc_0.start_buffer_0.start_buff.t3 VGND 0.060835f
C3921 tdc_0.start_buffer_0.start_buff.n20 VGND 0.449886f
C3922 tdc_0.start_buffer_0.start_buff.n21 VGND 0.114821f
C3923 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 VGND 0.09757f
C3924 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 VGND 0.030153f
C3925 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 VGND 0.265657f
C3926 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 VGND 0.039259f
C3927 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 VGND 0.012524f
C3928 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 VGND 0.027534f
C3929 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 VGND 0.039259f
C3930 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 VGND 0.012524f
C3931 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 VGND 0.027357f
C3932 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 VGND 0.008823f
C3933 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 VGND 0.039259f
C3934 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 VGND 0.012524f
C3935 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 VGND 0.027534f
C3936 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 VGND 0.039259f
C3937 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 VGND 0.012524f
C3938 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 VGND 0.027357f
C3939 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 VGND 0.008728f
C3940 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 VGND 0.135162f
C3941 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 VGND 0.046129f
C3942 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 VGND 0.046129f
C3943 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 VGND 0.054044f
C3944 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 VGND 0.046129f
C3945 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 VGND 0.046129f
C3946 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 VGND 0.0538f
C3947 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 VGND 0.495704f
C3948 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 VGND 0.119944f
C3949 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 VGND 0.025758f
C3950 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 VGND 0.025758f
C3951 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 VGND 0.055083f
C3952 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 VGND 0.008586f
C3953 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 VGND 0.008586f
C3954 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 VGND 0.01864f
C3955 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 VGND 0.221512f
C3956 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 VGND 0.09757f
C3957 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 VGND 0.030153f
C3958 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 VGND 0.234486f
C3959 tdc_0.vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n16 VGND 0.050613f
C3960 VDPWR.n0 VGND 0.078016f
C3961 VDPWR.t475 VGND 0.050452f
C3962 VDPWR.n1 VGND 0.114273f
C3963 VDPWR.n2 VGND 0.109479f
C3964 VDPWR.n3 VGND 0.109479f
C3965 VDPWR.t414 VGND 0.593337f
C3966 VDPWR.t474 VGND 0.015577f
C3967 VDPWR.n4 VGND 0.094938f
C3968 VDPWR.n5 VGND 0.074387f
C3969 VDPWR.n6 VGND 0.078004f
C3970 VDPWR.t1 VGND 0.050452f
C3971 VDPWR.n7 VGND 0.114273f
C3972 VDPWR.n8 VGND 0.109479f
C3973 VDPWR.n9 VGND 0.109479f
C3974 VDPWR.t165 VGND 0.590746f
C3975 VDPWR.t0 VGND 0.015509f
C3976 VDPWR.n10 VGND 0.094938f
C3977 VDPWR.n11 VGND 0.074387f
C3978 VDPWR.n12 VGND 0.046716f
C3979 VDPWR.t430 VGND 0.050473f
C3980 VDPWR.n13 VGND 0.052303f
C3981 VDPWR.n14 VGND 0.046716f
C3982 VDPWR.n15 VGND 0.030825f
C3983 VDPWR.n16 VGND 0.030825f
C3984 VDPWR.t429 VGND 0.460231f
C3985 VDPWR.n17 VGND 0.252266f
C3986 VDPWR.n18 VGND 0.030825f
C3987 VDPWR.n19 VGND 0.030825f
C3988 VDPWR.n20 VGND 0.046716f
C3989 VDPWR.n21 VGND 0.046716f
C3990 VDPWR.n22 VGND 0.05729f
C3991 VDPWR.t547 VGND 0.01345f
C3992 VDPWR.t278 VGND 0.01345f
C3993 VDPWR.n23 VGND 0.039254f
C3994 VDPWR.t380 VGND 0.049658f
C3995 VDPWR.n24 VGND 0.179043f
C3996 VDPWR.n25 VGND 0.07741f
C3997 VDPWR.n26 VGND 0.05729f
C3998 VDPWR.n27 VGND 0.036255f
C3999 VDPWR.n28 VGND 0.19772f
C4000 VDPWR.t548 VGND 0.168928f
C4001 VDPWR.n29 VGND 0.093512f
C4002 VDPWR.n30 VGND 0.07741f
C4003 VDPWR.t423 VGND 0.096114f
C4004 VDPWR.n31 VGND 0.064076f
C4005 VDPWR.t449 VGND 0.096114f
C4006 VDPWR.t438 VGND 0.189497f
C4007 VDPWR.n32 VGND 0.19772f
C4008 VDPWR.n33 VGND 0.05729f
C4009 VDPWR.t450 VGND 0.01345f
C4010 VDPWR.t424 VGND 0.01345f
C4011 VDPWR.n34 VGND 0.039254f
C4012 VDPWR.t439 VGND 0.049658f
C4013 VDPWR.n35 VGND 0.179043f
C4014 VDPWR.n36 VGND 0.046716f
C4015 VDPWR.t441 VGND 0.050473f
C4016 VDPWR.n37 VGND 0.052303f
C4017 VDPWR.n38 VGND 0.046716f
C4018 VDPWR.n39 VGND 0.030825f
C4019 VDPWR.n40 VGND 0.030825f
C4020 VDPWR.t137 VGND 0.460231f
C4021 VDPWR.n41 VGND 0.252266f
C4022 VDPWR.n42 VGND 0.030825f
C4023 VDPWR.n43 VGND 0.030825f
C4024 VDPWR.n44 VGND 0.048752f
C4025 VDPWR.n45 VGND 0.046716f
C4026 VDPWR.n46 VGND 0.05729f
C4027 VDPWR.t612 VGND 0.01345f
C4028 VDPWR.t610 VGND 0.01345f
C4029 VDPWR.n47 VGND 0.038685f
C4030 VDPWR.t485 VGND 0.049658f
C4031 VDPWR.n48 VGND 0.169321f
C4032 VDPWR.n49 VGND 0.07741f
C4033 VDPWR.n50 VGND 0.05729f
C4034 VDPWR.n51 VGND 0.036255f
C4035 VDPWR.n52 VGND 0.19772f
C4036 VDPWR.t84 VGND 0.168928f
C4037 VDPWR.n53 VGND 0.093512f
C4038 VDPWR.n54 VGND 0.07741f
C4039 VDPWR.t432 VGND 0.096114f
C4040 VDPWR.n55 VGND 0.064076f
C4041 VDPWR.t417 VGND 0.096114f
C4042 VDPWR.t446 VGND 0.189497f
C4043 VDPWR.n56 VGND 0.19772f
C4044 VDPWR.n57 VGND 0.057424f
C4045 VDPWR.t418 VGND 0.01345f
C4046 VDPWR.t433 VGND 0.01345f
C4047 VDPWR.n58 VGND 0.039254f
C4048 VDPWR.t447 VGND 0.049658f
C4049 VDPWR.n59 VGND 0.179043f
C4050 VDPWR.n60 VGND 0.036039f
C4051 VDPWR.n61 VGND 0.033541f
C4052 VDPWR.n62 VGND 0.093512f
C4053 VDPWR.n63 VGND 0.05729f
C4054 VDPWR.n64 VGND 0.036255f
C4055 VDPWR.n65 VGND 0.345136f
C4056 VDPWR.n66 VGND 0.345136f
C4057 VDPWR.t606 VGND 0.168928f
C4058 VDPWR.t611 VGND 0.096114f
C4059 VDPWR.t484 VGND 0.189497f
C4060 VDPWR.t609 VGND 0.096114f
C4061 VDPWR.n67 VGND 0.064076f
C4062 VDPWR.n68 VGND 0.093512f
C4063 VDPWR.n69 VGND 0.093512f
C4064 VDPWR.n70 VGND 0.033541f
C4065 VDPWR.n71 VGND 0.03641f
C4066 VDPWR.n72 VGND 0.043795f
C4067 VDPWR.n73 VGND 0.075724f
C4068 VDPWR.t138 VGND 0.050473f
C4069 VDPWR.n74 VGND 0.049038f
C4070 VDPWR.n75 VGND 0.093119f
C4071 VDPWR.n76 VGND 0.012244f
C4072 VDPWR.n77 VGND 0.060863f
C4073 VDPWR.n78 VGND 0.060863f
C4074 VDPWR.n79 VGND 0.340867f
C4075 VDPWR.n80 VGND 0.060863f
C4076 VDPWR.n81 VGND 0.060863f
C4077 VDPWR.n82 VGND 0.014025f
C4078 VDPWR.n83 VGND 0.093119f
C4079 VDPWR.n84 VGND 0.054058f
C4080 VDPWR.t440 VGND 0.020546f
C4081 VDPWR.t622 VGND 0.006632f
C4082 VDPWR.n85 VGND 0.020254f
C4083 VDPWR.t416 VGND 0.020267f
C4084 VDPWR.t445 VGND 0.021926f
C4085 VDPWR.n86 VGND 0.021512f
C4086 VDPWR.t431 VGND 0.021852f
C4087 VDPWR.n87 VGND 0.01497f
C4088 VDPWR.t624 VGND 0.006354f
C4089 VDPWR.t625 VGND 0.008155f
C4090 VDPWR.t632 VGND 0.008155f
C4091 VDPWR.n88 VGND 0.024443f
C4092 VDPWR.n89 VGND 0.150321f
C4093 VDPWR.n90 VGND 0.121093f
C4094 VDPWR.n91 VGND 0.147645f
C4095 VDPWR.n92 VGND 0.042318f
C4096 VDPWR.n93 VGND 0.036746f
C4097 VDPWR.n94 VGND 0.036039f
C4098 VDPWR.n95 VGND 0.033541f
C4099 VDPWR.n96 VGND 0.093512f
C4100 VDPWR.n97 VGND 0.05729f
C4101 VDPWR.n98 VGND 0.036255f
C4102 VDPWR.n99 VGND 0.345136f
C4103 VDPWR.n100 VGND 0.345136f
C4104 VDPWR.t115 VGND 0.168928f
C4105 VDPWR.t546 VGND 0.096114f
C4106 VDPWR.t379 VGND 0.189497f
C4107 VDPWR.t277 VGND 0.096114f
C4108 VDPWR.n101 VGND 0.064076f
C4109 VDPWR.n102 VGND 0.093512f
C4110 VDPWR.n103 VGND 0.093512f
C4111 VDPWR.n104 VGND 0.033541f
C4112 VDPWR.n105 VGND 0.03641f
C4113 VDPWR.n106 VGND 0.043795f
C4114 VDPWR.n107 VGND 0.073817f
C4115 VDPWR.t569 VGND 0.050473f
C4116 VDPWR.n108 VGND 0.049038f
C4117 VDPWR.n109 VGND 0.093119f
C4118 VDPWR.n110 VGND 0.014025f
C4119 VDPWR.n111 VGND 0.060863f
C4120 VDPWR.n112 VGND 0.060863f
C4121 VDPWR.n113 VGND 0.340867f
C4122 VDPWR.n114 VGND 0.060863f
C4123 VDPWR.n115 VGND 0.060863f
C4124 VDPWR.n116 VGND 0.014025f
C4125 VDPWR.n117 VGND 0.093119f
C4126 VDPWR.n118 VGND 0.055099f
C4127 VDPWR.t428 VGND 0.020546f
C4128 VDPWR.t626 VGND 0.006632f
C4129 VDPWR.n119 VGND 0.020264f
C4130 VDPWR.t448 VGND 0.020267f
C4131 VDPWR.t437 VGND 0.021926f
C4132 VDPWR.n120 VGND 0.021512f
C4133 VDPWR.t422 VGND 0.021852f
C4134 VDPWR.n121 VGND 0.01497f
C4135 VDPWR.t628 VGND 0.006354f
C4136 VDPWR.t630 VGND 0.008155f
C4137 VDPWR.t633 VGND 0.008155f
C4138 VDPWR.n122 VGND 0.024443f
C4139 VDPWR.n123 VGND 0.150321f
C4140 VDPWR.n124 VGND 0.120552f
C4141 VDPWR.n125 VGND 0.148176f
C4142 VDPWR.n126 VGND 0.029294f
C4143 VDPWR.n127 VGND 0.029946f
C4144 VDPWR.t166 VGND 0.050458f
C4145 VDPWR.n128 VGND 0.117901f
C4146 VDPWR.n129 VGND 0.236843f
C4147 VDPWR.n130 VGND 0.057418f
C4148 VDPWR.n131 VGND 0.041228f
C4149 VDPWR.n132 VGND 0.308156f
C4150 VDPWR.n133 VGND 0.025188f
C4151 VDPWR.n134 VGND 0.530186f
C4152 VDPWR.n135 VGND 0.099558f
C4153 VDPWR.n136 VGND 0.024488f
C4154 VDPWR.n137 VGND 0.109527f
C4155 VDPWR.n138 VGND 0.07145f
C4156 VDPWR.t415 VGND 0.050458f
C4157 VDPWR.n139 VGND 0.117901f
C4158 VDPWR.n140 VGND 0.116229f
C4159 VDPWR.n141 VGND 0.057418f
C4160 VDPWR.n142 VGND 0.041228f
C4161 VDPWR.n143 VGND 0.309542f
C4162 VDPWR.n144 VGND 0.025177f
C4163 VDPWR.n145 VGND 0.532041f
C4164 VDPWR.n146 VGND 0.099558f
C4165 VDPWR.n147 VGND 0.024488f
C4166 VDPWR.n148 VGND 0.109527f
C4167 VDPWR.n149 VGND 0.07145f
C4168 VDPWR.n150 VGND 0.10662f
C4169 VDPWR.n151 VGND 0.051039f
C4170 VDPWR.t608 VGND 0.050473f
C4171 VDPWR.n152 VGND 0.139191f
C4172 VDPWR.n153 VGND 0.22315f
C4173 VDPWR.t607 VGND 0.230116f
C4174 VDPWR.n154 VGND 0.030825f
C4175 VDPWR.n155 VGND 0.134279f
C4176 VDPWR.n156 VGND 0.019638f
C4177 VDPWR.n157 VGND 0.060869f
C4178 VDPWR.n158 VGND 0.060863f
C4179 VDPWR.n159 VGND 0.003488f
C4180 VDPWR.n160 VGND 0.072276f
C4181 VDPWR.n161 VGND 0.10078f
C4182 VDPWR.t532 VGND 0.050605f
C4183 VDPWR.n162 VGND 0.098879f
C4184 VDPWR.n163 VGND 0.075575f
C4185 VDPWR.n164 VGND 0.299591f
C4186 VDPWR.t531 VGND 0.28293f
C4187 VDPWR.t535 VGND 0.050605f
C4188 VDPWR.n165 VGND 0.01025f
C4189 VDPWR.n166 VGND 0.098879f
C4190 VDPWR.n167 VGND 0.060357f
C4191 VDPWR.t534 VGND 0.050468f
C4192 VDPWR.t427 VGND 0.050468f
C4193 VDPWR.n168 VGND 0.097282f
C4194 VDPWR.t627 VGND 0.015502f
C4195 VDPWR.t425 VGND 0.020899f
C4196 VDPWR.n169 VGND 0.023256f
C4197 VDPWR.n170 VGND 0.046665f
C4198 VDPWR.n171 VGND 0.078016f
C4199 VDPWR.t462 VGND 0.050452f
C4200 VDPWR.n172 VGND 0.114273f
C4201 VDPWR.n173 VGND 0.109479f
C4202 VDPWR.n174 VGND 0.109479f
C4203 VDPWR.t2 VGND 0.593337f
C4204 VDPWR.t461 VGND 0.015577f
C4205 VDPWR.n175 VGND 0.094938f
C4206 VDPWR.n176 VGND 0.074387f
C4207 VDPWR.n177 VGND 0.078004f
C4208 VDPWR.t17 VGND 0.050452f
C4209 VDPWR.n178 VGND 0.114273f
C4210 VDPWR.n179 VGND 0.109479f
C4211 VDPWR.n180 VGND 0.109479f
C4212 VDPWR.t76 VGND 0.590746f
C4213 VDPWR.t16 VGND 0.015509f
C4214 VDPWR.n181 VGND 0.094938f
C4215 VDPWR.n182 VGND 0.074387f
C4216 VDPWR.n183 VGND 0.046716f
C4217 VDPWR.t151 VGND 0.050473f
C4218 VDPWR.n184 VGND 0.052303f
C4219 VDPWR.n185 VGND 0.046716f
C4220 VDPWR.n186 VGND 0.030825f
C4221 VDPWR.n187 VGND 0.030825f
C4222 VDPWR.t150 VGND 0.460231f
C4223 VDPWR.n188 VGND 0.252266f
C4224 VDPWR.n189 VGND 0.030825f
C4225 VDPWR.n190 VGND 0.030825f
C4226 VDPWR.n191 VGND 0.046716f
C4227 VDPWR.n192 VGND 0.046716f
C4228 VDPWR.n193 VGND 0.05729f
C4229 VDPWR.t593 VGND 0.01345f
C4230 VDPWR.t342 VGND 0.01345f
C4231 VDPWR.n194 VGND 0.039254f
C4232 VDPWR.t340 VGND 0.049658f
C4233 VDPWR.n195 VGND 0.179043f
C4234 VDPWR.n196 VGND 0.07741f
C4235 VDPWR.n197 VGND 0.05729f
C4236 VDPWR.n198 VGND 0.036255f
C4237 VDPWR.n199 VGND 0.19772f
C4238 VDPWR.t39 VGND 0.168928f
C4239 VDPWR.n200 VGND 0.093512f
C4240 VDPWR.n201 VGND 0.07741f
C4241 VDPWR.t148 VGND 0.096114f
C4242 VDPWR.n202 VGND 0.064076f
C4243 VDPWR.t221 VGND 0.096114f
C4244 VDPWR.t477 VGND 0.189497f
C4245 VDPWR.n203 VGND 0.19772f
C4246 VDPWR.n204 VGND 0.05729f
C4247 VDPWR.t222 VGND 0.01345f
C4248 VDPWR.t149 VGND 0.01345f
C4249 VDPWR.n205 VGND 0.039254f
C4250 VDPWR.t478 VGND 0.049658f
C4251 VDPWR.n206 VGND 0.179043f
C4252 VDPWR.n207 VGND 0.046716f
C4253 VDPWR.t533 VGND 0.050473f
C4254 VDPWR.n208 VGND 0.052303f
C4255 VDPWR.n209 VGND 0.046716f
C4256 VDPWR.n210 VGND 0.030825f
C4257 VDPWR.n211 VGND 0.030825f
C4258 VDPWR.t527 VGND 0.460231f
C4259 VDPWR.n212 VGND 0.252266f
C4260 VDPWR.n213 VGND 0.030825f
C4261 VDPWR.n214 VGND 0.030825f
C4262 VDPWR.n215 VGND 0.046716f
C4263 VDPWR.n216 VGND 0.046716f
C4264 VDPWR.n217 VGND 0.05729f
C4265 VDPWR.t95 VGND 0.01345f
C4266 VDPWR.t406 VGND 0.01345f
C4267 VDPWR.n218 VGND 0.039254f
C4268 VDPWR.t503 VGND 0.049658f
C4269 VDPWR.n219 VGND 0.179043f
C4270 VDPWR.n220 VGND 0.07741f
C4271 VDPWR.n221 VGND 0.05729f
C4272 VDPWR.n222 VGND 0.036255f
C4273 VDPWR.n223 VGND 0.19772f
C4274 VDPWR.t61 VGND 0.168928f
C4275 VDPWR.n224 VGND 0.093512f
C4276 VDPWR.n225 VGND 0.07741f
C4277 VDPWR.t357 VGND 0.096114f
C4278 VDPWR.n226 VGND 0.064076f
C4279 VDPWR.t265 VGND 0.096114f
C4280 VDPWR.t575 VGND 0.189497f
C4281 VDPWR.n227 VGND 0.19772f
C4282 VDPWR.n228 VGND 0.05729f
C4283 VDPWR.t266 VGND 0.01345f
C4284 VDPWR.t358 VGND 0.01345f
C4285 VDPWR.n229 VGND 0.039254f
C4286 VDPWR.t576 VGND 0.049658f
C4287 VDPWR.n230 VGND 0.179043f
C4288 VDPWR.n231 VGND 0.046716f
C4289 VDPWR.t306 VGND 0.050473f
C4290 VDPWR.n232 VGND 0.052303f
C4291 VDPWR.n233 VGND 0.046716f
C4292 VDPWR.n234 VGND 0.030825f
C4293 VDPWR.n235 VGND 0.030825f
C4294 VDPWR.t305 VGND 0.460231f
C4295 VDPWR.n236 VGND 0.252266f
C4296 VDPWR.n237 VGND 0.030825f
C4297 VDPWR.n238 VGND 0.030825f
C4298 VDPWR.n239 VGND 0.046716f
C4299 VDPWR.n240 VGND 0.046716f
C4300 VDPWR.n241 VGND 0.05729f
C4301 VDPWR.t259 VGND 0.01345f
C4302 VDPWR.t257 VGND 0.01345f
C4303 VDPWR.n242 VGND 0.039254f
C4304 VDPWR.t327 VGND 0.049658f
C4305 VDPWR.n243 VGND 0.179043f
C4306 VDPWR.n244 VGND 0.07741f
C4307 VDPWR.n245 VGND 0.05729f
C4308 VDPWR.n246 VGND 0.036255f
C4309 VDPWR.n247 VGND 0.19772f
C4310 VDPWR.t42 VGND 0.168928f
C4311 VDPWR.n248 VGND 0.093512f
C4312 VDPWR.n249 VGND 0.07741f
C4313 VDPWR.t51 VGND 0.096114f
C4314 VDPWR.n250 VGND 0.064076f
C4315 VDPWR.t78 VGND 0.096114f
C4316 VDPWR.t80 VGND 0.189497f
C4317 VDPWR.n251 VGND 0.19772f
C4318 VDPWR.n252 VGND 0.05729f
C4319 VDPWR.t79 VGND 0.01345f
C4320 VDPWR.t52 VGND 0.01345f
C4321 VDPWR.n253 VGND 0.039254f
C4322 VDPWR.t81 VGND 0.049658f
C4323 VDPWR.n254 VGND 0.179043f
C4324 VDPWR.n255 VGND 0.046716f
C4325 VDPWR.t184 VGND 0.050473f
C4326 VDPWR.n256 VGND 0.052303f
C4327 VDPWR.n257 VGND 0.046716f
C4328 VDPWR.n258 VGND 0.030825f
C4329 VDPWR.n259 VGND 0.030825f
C4330 VDPWR.t74 VGND 0.460231f
C4331 VDPWR.n260 VGND 0.252266f
C4332 VDPWR.n261 VGND 0.030825f
C4333 VDPWR.n262 VGND 0.030825f
C4334 VDPWR.n263 VGND 0.046716f
C4335 VDPWR.n264 VGND 0.046716f
C4336 VDPWR.n265 VGND 0.05729f
C4337 VDPWR.t245 VGND 0.01345f
C4338 VDPWR.t356 VGND 0.01345f
C4339 VDPWR.n266 VGND 0.039254f
C4340 VDPWR.t354 VGND 0.049658f
C4341 VDPWR.n267 VGND 0.179043f
C4342 VDPWR.n268 VGND 0.07741f
C4343 VDPWR.n269 VGND 0.05729f
C4344 VDPWR.n270 VGND 0.036255f
C4345 VDPWR.n271 VGND 0.19772f
C4346 VDPWR.t473 VGND 0.168928f
C4347 VDPWR.n272 VGND 0.093512f
C4348 VDPWR.n273 VGND 0.07741f
C4349 VDPWR.t274 VGND 0.096114f
C4350 VDPWR.n274 VGND 0.064076f
C4351 VDPWR.t554 VGND 0.096114f
C4352 VDPWR.t552 VGND 0.189497f
C4353 VDPWR.n275 VGND 0.19772f
C4354 VDPWR.n276 VGND 0.05729f
C4355 VDPWR.t555 VGND 0.01345f
C4356 VDPWR.t275 VGND 0.01345f
C4357 VDPWR.n277 VGND 0.039254f
C4358 VDPWR.t553 VGND 0.049658f
C4359 VDPWR.n278 VGND 0.179043f
C4360 VDPWR.n279 VGND 0.046716f
C4361 VDPWR.t122 VGND 0.050473f
C4362 VDPWR.n280 VGND 0.052303f
C4363 VDPWR.n281 VGND 0.046716f
C4364 VDPWR.n282 VGND 0.030825f
C4365 VDPWR.n283 VGND 0.030825f
C4366 VDPWR.t70 VGND 0.460231f
C4367 VDPWR.n284 VGND 0.252266f
C4368 VDPWR.n285 VGND 0.030825f
C4369 VDPWR.n286 VGND 0.030825f
C4370 VDPWR.n287 VGND 0.046716f
C4371 VDPWR.n288 VGND 0.046716f
C4372 VDPWR.n289 VGND 0.05729f
C4373 VDPWR.t203 VGND 0.01345f
C4374 VDPWR.t413 VGND 0.01345f
C4375 VDPWR.n290 VGND 0.039254f
C4376 VDPWR.t205 VGND 0.049658f
C4377 VDPWR.n291 VGND 0.179043f
C4378 VDPWR.n292 VGND 0.07741f
C4379 VDPWR.n293 VGND 0.05729f
C4380 VDPWR.n294 VGND 0.036255f
C4381 VDPWR.n295 VGND 0.19772f
C4382 VDPWR.t14 VGND 0.168928f
C4383 VDPWR.n296 VGND 0.093512f
C4384 VDPWR.n297 VGND 0.07741f
C4385 VDPWR.t514 VGND 0.096114f
C4386 VDPWR.n298 VGND 0.064076f
C4387 VDPWR.t123 VGND 0.096114f
C4388 VDPWR.t120 VGND 0.189497f
C4389 VDPWR.n299 VGND 0.19772f
C4390 VDPWR.n300 VGND 0.05729f
C4391 VDPWR.t124 VGND 0.01345f
C4392 VDPWR.t515 VGND 0.01345f
C4393 VDPWR.n301 VGND 0.039254f
C4394 VDPWR.t121 VGND 0.049658f
C4395 VDPWR.n302 VGND 0.179043f
C4396 VDPWR.n303 VGND 0.046716f
C4397 VDPWR.t452 VGND 0.050473f
C4398 VDPWR.n304 VGND 0.052303f
C4399 VDPWR.n305 VGND 0.046716f
C4400 VDPWR.n306 VGND 0.030825f
C4401 VDPWR.n307 VGND 0.030825f
C4402 VDPWR.t254 VGND 0.460231f
C4403 VDPWR.n308 VGND 0.252266f
C4404 VDPWR.n309 VGND 0.030825f
C4405 VDPWR.n310 VGND 0.030825f
C4406 VDPWR.n311 VGND 0.046716f
C4407 VDPWR.n312 VGND 0.046716f
C4408 VDPWR.n313 VGND 0.05729f
C4409 VDPWR.t509 VGND 0.01345f
C4410 VDPWR.t352 VGND 0.01345f
C4411 VDPWR.n314 VGND 0.039254f
C4412 VDPWR.t243 VGND 0.049658f
C4413 VDPWR.n315 VGND 0.179043f
C4414 VDPWR.n316 VGND 0.07741f
C4415 VDPWR.n317 VGND 0.05729f
C4416 VDPWR.n318 VGND 0.036255f
C4417 VDPWR.n319 VGND 0.19772f
C4418 VDPWR.t83 VGND 0.168928f
C4419 VDPWR.n320 VGND 0.093512f
C4420 VDPWR.n321 VGND 0.07741f
C4421 VDPWR.t435 VGND 0.096114f
C4422 VDPWR.n322 VGND 0.064076f
C4423 VDPWR.t420 VGND 0.096114f
C4424 VDPWR.t443 VGND 0.189497f
C4425 VDPWR.n323 VGND 0.19772f
C4426 VDPWR.n324 VGND 0.057424f
C4427 VDPWR.t421 VGND 0.01345f
C4428 VDPWR.t436 VGND 0.01345f
C4429 VDPWR.n325 VGND 0.039254f
C4430 VDPWR.t444 VGND 0.049658f
C4431 VDPWR.n326 VGND 0.179043f
C4432 VDPWR.n327 VGND 0.036039f
C4433 VDPWR.n328 VGND 0.033541f
C4434 VDPWR.n329 VGND 0.093512f
C4435 VDPWR.n330 VGND 0.05729f
C4436 VDPWR.n331 VGND 0.036255f
C4437 VDPWR.n332 VGND 0.345136f
C4438 VDPWR.n333 VGND 0.345136f
C4439 VDPWR.t100 VGND 0.168928f
C4440 VDPWR.t508 VGND 0.096114f
C4441 VDPWR.t242 VGND 0.189497f
C4442 VDPWR.t351 VGND 0.096114f
C4443 VDPWR.n334 VGND 0.064076f
C4444 VDPWR.n335 VGND 0.093512f
C4445 VDPWR.n336 VGND 0.093512f
C4446 VDPWR.n337 VGND 0.033541f
C4447 VDPWR.n338 VGND 0.03641f
C4448 VDPWR.n339 VGND 0.043795f
C4449 VDPWR.n340 VGND 0.073817f
C4450 VDPWR.t255 VGND 0.050473f
C4451 VDPWR.n341 VGND 0.049038f
C4452 VDPWR.n342 VGND 0.093119f
C4453 VDPWR.n343 VGND 0.014025f
C4454 VDPWR.n344 VGND 0.060863f
C4455 VDPWR.n345 VGND 0.060863f
C4456 VDPWR.n346 VGND 0.340867f
C4457 VDPWR.n347 VGND 0.060863f
C4458 VDPWR.n348 VGND 0.060863f
C4459 VDPWR.n349 VGND 0.014025f
C4460 VDPWR.n350 VGND 0.093119f
C4461 VDPWR.n351 VGND 0.053737f
C4462 VDPWR.t451 VGND 0.020546f
C4463 VDPWR.t621 VGND 0.006632f
C4464 VDPWR.n352 VGND 0.020251f
C4465 VDPWR.t419 VGND 0.020267f
C4466 VDPWR.t442 VGND 0.021926f
C4467 VDPWR.n353 VGND 0.021512f
C4468 VDPWR.t434 VGND 0.021852f
C4469 VDPWR.n354 VGND 0.01497f
C4470 VDPWR.t631 VGND 0.006354f
C4471 VDPWR.t623 VGND 0.008155f
C4472 VDPWR.t629 VGND 0.008155f
C4473 VDPWR.n355 VGND 0.024443f
C4474 VDPWR.n356 VGND 0.150321f
C4475 VDPWR.n357 VGND 0.121256f
C4476 VDPWR.n358 VGND 0.147486f
C4477 VDPWR.n359 VGND 0.042361f
C4478 VDPWR.n360 VGND 0.036746f
C4479 VDPWR.n361 VGND 0.036039f
C4480 VDPWR.n362 VGND 0.033541f
C4481 VDPWR.n363 VGND 0.093512f
C4482 VDPWR.n364 VGND 0.05729f
C4483 VDPWR.n365 VGND 0.036255f
C4484 VDPWR.n366 VGND 0.345136f
C4485 VDPWR.n367 VGND 0.345136f
C4486 VDPWR.t579 VGND 0.168928f
C4487 VDPWR.t202 VGND 0.096114f
C4488 VDPWR.t204 VGND 0.189497f
C4489 VDPWR.t412 VGND 0.096114f
C4490 VDPWR.n368 VGND 0.064076f
C4491 VDPWR.n369 VGND 0.093512f
C4492 VDPWR.n370 VGND 0.093512f
C4493 VDPWR.n371 VGND 0.033541f
C4494 VDPWR.n372 VGND 0.03641f
C4495 VDPWR.n373 VGND 0.043795f
C4496 VDPWR.n374 VGND 0.073817f
C4497 VDPWR.t71 VGND 0.050473f
C4498 VDPWR.n375 VGND 0.049038f
C4499 VDPWR.n376 VGND 0.093119f
C4500 VDPWR.n377 VGND 0.014025f
C4501 VDPWR.n378 VGND 0.060863f
C4502 VDPWR.n379 VGND 0.060863f
C4503 VDPWR.n380 VGND 0.340867f
C4504 VDPWR.n381 VGND 0.060863f
C4505 VDPWR.n382 VGND 0.060863f
C4506 VDPWR.n383 VGND 0.014025f
C4507 VDPWR.n384 VGND 0.093119f
C4508 VDPWR.n385 VGND 0.082788f
C4509 VDPWR.n386 VGND 0.036746f
C4510 VDPWR.n387 VGND 0.036039f
C4511 VDPWR.n388 VGND 0.033541f
C4512 VDPWR.n389 VGND 0.093512f
C4513 VDPWR.n390 VGND 0.05729f
C4514 VDPWR.n391 VGND 0.036255f
C4515 VDPWR.n392 VGND 0.345136f
C4516 VDPWR.n393 VGND 0.345136f
C4517 VDPWR.t125 VGND 0.168928f
C4518 VDPWR.t244 VGND 0.096114f
C4519 VDPWR.t353 VGND 0.189497f
C4520 VDPWR.t355 VGND 0.096114f
C4521 VDPWR.n394 VGND 0.064076f
C4522 VDPWR.n395 VGND 0.093512f
C4523 VDPWR.n396 VGND 0.093512f
C4524 VDPWR.n397 VGND 0.033541f
C4525 VDPWR.n398 VGND 0.03641f
C4526 VDPWR.n399 VGND 0.043795f
C4527 VDPWR.n400 VGND 0.073817f
C4528 VDPWR.t75 VGND 0.050473f
C4529 VDPWR.n401 VGND 0.049038f
C4530 VDPWR.n402 VGND 0.093119f
C4531 VDPWR.n403 VGND 0.014025f
C4532 VDPWR.n404 VGND 0.060863f
C4533 VDPWR.n405 VGND 0.060863f
C4534 VDPWR.n406 VGND 0.340867f
C4535 VDPWR.n407 VGND 0.060863f
C4536 VDPWR.n408 VGND 0.060863f
C4537 VDPWR.n409 VGND 0.014025f
C4538 VDPWR.n410 VGND 0.093119f
C4539 VDPWR.n411 VGND 0.082788f
C4540 VDPWR.n412 VGND 0.036746f
C4541 VDPWR.n413 VGND 0.036039f
C4542 VDPWR.n414 VGND 0.033541f
C4543 VDPWR.n415 VGND 0.093512f
C4544 VDPWR.n416 VGND 0.05729f
C4545 VDPWR.n417 VGND 0.036255f
C4546 VDPWR.n418 VGND 0.345136f
C4547 VDPWR.n419 VGND 0.345136f
C4548 VDPWR.t289 VGND 0.168928f
C4549 VDPWR.t258 VGND 0.096114f
C4550 VDPWR.t326 VGND 0.189497f
C4551 VDPWR.t256 VGND 0.096114f
C4552 VDPWR.n420 VGND 0.064076f
C4553 VDPWR.n421 VGND 0.093512f
C4554 VDPWR.n422 VGND 0.093512f
C4555 VDPWR.n423 VGND 0.033541f
C4556 VDPWR.n424 VGND 0.03641f
C4557 VDPWR.n425 VGND 0.043795f
C4558 VDPWR.n426 VGND 0.073817f
C4559 VDPWR.t549 VGND 0.050473f
C4560 VDPWR.n427 VGND 0.049038f
C4561 VDPWR.n428 VGND 0.093119f
C4562 VDPWR.n429 VGND 0.014025f
C4563 VDPWR.n430 VGND 0.060863f
C4564 VDPWR.n431 VGND 0.060863f
C4565 VDPWR.n432 VGND 0.340867f
C4566 VDPWR.n433 VGND 0.060863f
C4567 VDPWR.n434 VGND 0.060863f
C4568 VDPWR.n435 VGND 0.014025f
C4569 VDPWR.n436 VGND 0.093119f
C4570 VDPWR.n437 VGND 0.082788f
C4571 VDPWR.n438 VGND 0.036746f
C4572 VDPWR.n439 VGND 0.036039f
C4573 VDPWR.n440 VGND 0.033541f
C4574 VDPWR.n441 VGND 0.093512f
C4575 VDPWR.n442 VGND 0.05729f
C4576 VDPWR.n443 VGND 0.036255f
C4577 VDPWR.n444 VGND 0.345136f
C4578 VDPWR.n445 VGND 0.345136f
C4579 VDPWR.t516 VGND 0.168928f
C4580 VDPWR.t94 VGND 0.096114f
C4581 VDPWR.t502 VGND 0.189497f
C4582 VDPWR.t405 VGND 0.096114f
C4583 VDPWR.n446 VGND 0.064076f
C4584 VDPWR.n447 VGND 0.093512f
C4585 VDPWR.n448 VGND 0.093512f
C4586 VDPWR.n449 VGND 0.033541f
C4587 VDPWR.n450 VGND 0.03641f
C4588 VDPWR.n451 VGND 0.043795f
C4589 VDPWR.n452 VGND 0.073817f
C4590 VDPWR.t528 VGND 0.050473f
C4591 VDPWR.n453 VGND 0.049038f
C4592 VDPWR.n454 VGND 0.093119f
C4593 VDPWR.n455 VGND 0.014025f
C4594 VDPWR.n456 VGND 0.060863f
C4595 VDPWR.n457 VGND 0.060863f
C4596 VDPWR.n458 VGND 0.340867f
C4597 VDPWR.n459 VGND 0.060863f
C4598 VDPWR.n460 VGND 0.060863f
C4599 VDPWR.n461 VGND 0.014025f
C4600 VDPWR.n462 VGND 0.093119f
C4601 VDPWR.n463 VGND 0.082788f
C4602 VDPWR.n464 VGND 0.036746f
C4603 VDPWR.n465 VGND 0.036039f
C4604 VDPWR.n466 VGND 0.033541f
C4605 VDPWR.n467 VGND 0.093512f
C4606 VDPWR.n468 VGND 0.05729f
C4607 VDPWR.n469 VGND 0.036255f
C4608 VDPWR.n470 VGND 0.345136f
C4609 VDPWR.n471 VGND 0.345136f
C4610 VDPWR.t233 VGND 0.168928f
C4611 VDPWR.t592 VGND 0.096114f
C4612 VDPWR.t339 VGND 0.189497f
C4613 VDPWR.t341 VGND 0.096114f
C4614 VDPWR.n472 VGND 0.064076f
C4615 VDPWR.n473 VGND 0.093512f
C4616 VDPWR.n474 VGND 0.093512f
C4617 VDPWR.n475 VGND 0.033541f
C4618 VDPWR.n476 VGND 0.03641f
C4619 VDPWR.n477 VGND 0.043795f
C4620 VDPWR.n478 VGND 0.073817f
C4621 VDPWR.t300 VGND 0.050473f
C4622 VDPWR.n479 VGND 0.049038f
C4623 VDPWR.n480 VGND 0.093119f
C4624 VDPWR.n481 VGND 0.014025f
C4625 VDPWR.n482 VGND 0.060863f
C4626 VDPWR.n483 VGND 0.060863f
C4627 VDPWR.n484 VGND 0.340867f
C4628 VDPWR.n485 VGND 0.060863f
C4629 VDPWR.n486 VGND 0.060863f
C4630 VDPWR.n487 VGND 0.014025f
C4631 VDPWR.n488 VGND 0.093119f
C4632 VDPWR.n489 VGND 0.067907f
C4633 VDPWR.n490 VGND 0.04606f
C4634 VDPWR.t77 VGND 0.050458f
C4635 VDPWR.n491 VGND 0.117901f
C4636 VDPWR.n492 VGND 0.219321f
C4637 VDPWR.n493 VGND 0.057418f
C4638 VDPWR.n494 VGND 0.041228f
C4639 VDPWR.n495 VGND 0.308156f
C4640 VDPWR.n496 VGND 0.025188f
C4641 VDPWR.n497 VGND 0.530186f
C4642 VDPWR.n498 VGND 0.099558f
C4643 VDPWR.n499 VGND 0.024488f
C4644 VDPWR.n500 VGND 0.109527f
C4645 VDPWR.n501 VGND 0.07145f
C4646 VDPWR.t3 VGND 0.050458f
C4647 VDPWR.n502 VGND 0.117901f
C4648 VDPWR.n503 VGND 0.116229f
C4649 VDPWR.n504 VGND 0.057418f
C4650 VDPWR.n505 VGND 0.041228f
C4651 VDPWR.n506 VGND 0.309542f
C4652 VDPWR.n507 VGND 0.025177f
C4653 VDPWR.n508 VGND 0.532041f
C4654 VDPWR.n509 VGND 0.099558f
C4655 VDPWR.n510 VGND 0.024488f
C4656 VDPWR.n511 VGND 0.109527f
C4657 VDPWR.n512 VGND 0.07145f
C4658 VDPWR.n513 VGND 0.10662f
C4659 VDPWR.n514 VGND 0.051039f
C4660 VDPWR.t153 VGND 0.050473f
C4661 VDPWR.n515 VGND 0.139191f
C4662 VDPWR.n516 VGND 0.22315f
C4663 VDPWR.t152 VGND 0.230116f
C4664 VDPWR.n517 VGND 0.030825f
C4665 VDPWR.n518 VGND 0.134279f
C4666 VDPWR.n519 VGND 0.019638f
C4667 VDPWR.n520 VGND 0.060869f
C4668 VDPWR.n521 VGND 0.060863f
C4669 VDPWR.n522 VGND 0.003488f
C4670 VDPWR.n523 VGND 0.072276f
C4671 VDPWR.n524 VGND 0.095418f
C4672 VDPWR.n525 VGND 0.079082f
C4673 VDPWR.n526 VGND 0.042364f
C4674 VDPWR.n527 VGND 0.04794f
C4675 VDPWR.n528 VGND 0.032123f
C4676 VDPWR.t426 VGND 0.28293f
C4677 VDPWR.n529 VGND 0.161177f
C4678 VDPWR.n530 VGND 0.019706f
C4679 VDPWR.n531 VGND 0.299591f
C4680 VDPWR.n532 VGND 0.075575f
C4681 VDPWR.n533 VGND 0.013876f
C4682 VDPWR.n534 VGND 0.097282f
C4683 VDPWR.n535 VGND 1.11337f
C4684 VDPWR.t291 VGND 0.050838f
C4685 VDPWR.t319 VGND 0.050471f
C4686 VDPWR.n536 VGND 0.187611f
C4687 VDPWR.t119 VGND 0.050471f
C4688 VDPWR.n537 VGND 0.099429f
C4689 VDPWR.t145 VGND 0.050471f
C4690 VDPWR.n538 VGND 0.094949f
C4691 VDPWR.n539 VGND 0.062139f
C4692 VDPWR.n540 VGND 0.037271f
C4693 VDPWR.t216 VGND 0.050838f
C4694 VDPWR.t407 VGND 0.050471f
C4695 VDPWR.n541 VGND 0.187611f
C4696 VDPWR.t343 VGND 0.050471f
C4697 VDPWR.n542 VGND 0.099429f
C4698 VDPWR.t186 VGND 0.050471f
C4699 VDPWR.n543 VGND 0.094949f
C4700 VDPWR.n544 VGND 0.062139f
C4701 VDPWR.n545 VGND 0.037271f
C4702 VDPWR.t479 VGND 0.050838f
C4703 VDPWR.t170 VGND 0.050471f
C4704 VDPWR.n546 VGND 0.187611f
C4705 VDPWR.t334 VGND 0.050471f
C4706 VDPWR.n547 VGND 0.099429f
C4707 VDPWR.t285 VGND 0.050471f
C4708 VDPWR.n548 VGND 0.094949f
C4709 VDPWR.n549 VGND 0.062139f
C4710 VDPWR.n550 VGND 0.037271f
C4711 VDPWR.t486 VGND 0.050838f
C4712 VDPWR.t157 VGND 0.050471f
C4713 VDPWR.n551 VGND 0.187611f
C4714 VDPWR.t199 VGND 0.050471f
C4715 VDPWR.n552 VGND 0.099429f
C4716 VDPWR.t493 VGND 0.050471f
C4717 VDPWR.n553 VGND 0.094949f
C4718 VDPWR.n554 VGND 0.062139f
C4719 VDPWR.n555 VGND 0.037271f
C4720 VDPWR.t188 VGND 0.050838f
C4721 VDPWR.t583 VGND 0.050471f
C4722 VDPWR.n556 VGND 0.187611f
C4723 VDPWR.t276 VGND 0.050471f
C4724 VDPWR.n557 VGND 0.099429f
C4725 VDPWR.t381 VGND 0.050471f
C4726 VDPWR.n558 VGND 0.094949f
C4727 VDPWR.n559 VGND 0.062139f
C4728 VDPWR.n560 VGND 0.037271f
C4729 VDPWR.t286 VGND 0.050838f
C4730 VDPWR.t348 VGND 0.050471f
C4731 VDPWR.n561 VGND 0.187611f
C4732 VDPWR.t226 VGND 0.050471f
C4733 VDPWR.n562 VGND 0.099429f
C4734 VDPWR.t215 VGND 0.050471f
C4735 VDPWR.n563 VGND 0.094949f
C4736 VDPWR.n564 VGND 0.062139f
C4737 VDPWR.n565 VGND 0.037271f
C4738 VDPWR.t396 VGND 0.050838f
C4739 VDPWR.t293 VGND 0.050471f
C4740 VDPWR.n566 VGND 0.187611f
C4741 VDPWR.t99 VGND 0.050471f
C4742 VDPWR.n567 VGND 0.099429f
C4743 VDPWR.t292 VGND 0.050471f
C4744 VDPWR.n568 VGND 0.094949f
C4745 VDPWR.n569 VGND 0.062139f
C4746 VDPWR.n570 VGND 0.037271f
C4747 VDPWR.t283 VGND 0.050838f
C4748 VDPWR.t104 VGND 0.050471f
C4749 VDPWR.n571 VGND 0.187611f
C4750 VDPWR.t580 VGND 0.050471f
C4751 VDPWR.n572 VGND 0.099429f
C4752 VDPWR.t114 VGND 0.050471f
C4753 VDPWR.n573 VGND 0.094949f
C4754 VDPWR.n574 VGND 0.268877f
C4755 VDPWR.n575 VGND 0.037271f
C4756 VDPWR.n576 VGND 0.306591f
C4757 VDPWR.n577 VGND 0.121863f
C4758 VDPWR.t103 VGND 0.66253f
C4759 VDPWR.n578 VGND 0.155747f
C4760 VDPWR.n579 VGND 0.371223f
C4761 VDPWR.n580 VGND 0.39542f
C4762 VDPWR.n581 VGND 0.041768f
C4763 VDPWR.n582 VGND 0.036489f
C4764 VDPWR.n583 VGND 0.041768f
C4765 VDPWR.n584 VGND 0.073918f
C4766 VDPWR.n585 VGND 0.046407f
C4767 VDPWR.n586 VGND 0.006601f
C4768 VDPWR.n587 VGND 0.503555f
C4769 VDPWR.n588 VGND 0.078633f
C4770 VDPWR.n589 VGND 0.078633f
C4771 VDPWR.n590 VGND 0.065925f
C4772 VDPWR.n591 VGND 0.107512f
C4773 VDPWR.n592 VGND 0.202734f
C4774 VDPWR.n593 VGND 0.149751f
C4775 VDPWR.n594 VGND 0.121863f
C4776 VDPWR.t98 VGND 0.66253f
C4777 VDPWR.n595 VGND 0.155747f
C4778 VDPWR.n596 VGND 0.371223f
C4779 VDPWR.n597 VGND 0.39542f
C4780 VDPWR.n598 VGND 0.041768f
C4781 VDPWR.n599 VGND 0.036489f
C4782 VDPWR.n600 VGND 0.041768f
C4783 VDPWR.n601 VGND 0.073918f
C4784 VDPWR.n602 VGND 0.046407f
C4785 VDPWR.n603 VGND 0.006601f
C4786 VDPWR.n604 VGND 0.503555f
C4787 VDPWR.n605 VGND 0.078633f
C4788 VDPWR.n606 VGND 0.078633f
C4789 VDPWR.n607 VGND 0.065925f
C4790 VDPWR.n608 VGND 0.107512f
C4791 VDPWR.n609 VGND 0.202734f
C4792 VDPWR.n610 VGND 0.149751f
C4793 VDPWR.n611 VGND 0.121863f
C4794 VDPWR.t214 VGND 0.66253f
C4795 VDPWR.n612 VGND 0.155747f
C4796 VDPWR.n613 VGND 0.371223f
C4797 VDPWR.n614 VGND 0.39542f
C4798 VDPWR.n615 VGND 0.041768f
C4799 VDPWR.n616 VGND 0.036489f
C4800 VDPWR.n617 VGND 0.041768f
C4801 VDPWR.n618 VGND 0.073918f
C4802 VDPWR.n619 VGND 0.046407f
C4803 VDPWR.n620 VGND 0.006601f
C4804 VDPWR.n621 VGND 0.503555f
C4805 VDPWR.n622 VGND 0.078633f
C4806 VDPWR.n623 VGND 0.078633f
C4807 VDPWR.n624 VGND 0.065925f
C4808 VDPWR.n625 VGND 0.107512f
C4809 VDPWR.n626 VGND 0.202734f
C4810 VDPWR.n627 VGND 0.149751f
C4811 VDPWR.n628 VGND 0.121863f
C4812 VDPWR.t187 VGND 0.66253f
C4813 VDPWR.n629 VGND 0.155747f
C4814 VDPWR.n630 VGND 0.371223f
C4815 VDPWR.n631 VGND 0.39542f
C4816 VDPWR.n632 VGND 0.041768f
C4817 VDPWR.n633 VGND 0.036489f
C4818 VDPWR.n634 VGND 0.041768f
C4819 VDPWR.n635 VGND 0.073918f
C4820 VDPWR.n636 VGND 0.046407f
C4821 VDPWR.n637 VGND 0.006601f
C4822 VDPWR.n638 VGND 0.503555f
C4823 VDPWR.n639 VGND 0.078633f
C4824 VDPWR.n640 VGND 0.078633f
C4825 VDPWR.n641 VGND 0.065925f
C4826 VDPWR.n642 VGND 0.107512f
C4827 VDPWR.n643 VGND 0.202734f
C4828 VDPWR.n644 VGND 0.149751f
C4829 VDPWR.n645 VGND 0.121863f
C4830 VDPWR.t156 VGND 0.66253f
C4831 VDPWR.n646 VGND 0.155747f
C4832 VDPWR.n647 VGND 0.371223f
C4833 VDPWR.n648 VGND 0.39542f
C4834 VDPWR.n649 VGND 0.041768f
C4835 VDPWR.n650 VGND 0.036489f
C4836 VDPWR.n651 VGND 0.041768f
C4837 VDPWR.n652 VGND 0.073918f
C4838 VDPWR.n653 VGND 0.046407f
C4839 VDPWR.n654 VGND 0.006601f
C4840 VDPWR.n655 VGND 0.503555f
C4841 VDPWR.n656 VGND 0.078633f
C4842 VDPWR.n657 VGND 0.078633f
C4843 VDPWR.n658 VGND 0.065925f
C4844 VDPWR.n659 VGND 0.107512f
C4845 VDPWR.n660 VGND 0.202734f
C4846 VDPWR.n661 VGND 0.149751f
C4847 VDPWR.n662 VGND 0.121863f
C4848 VDPWR.t169 VGND 0.66253f
C4849 VDPWR.n663 VGND 0.155747f
C4850 VDPWR.n664 VGND 0.371223f
C4851 VDPWR.n665 VGND 0.39542f
C4852 VDPWR.n666 VGND 0.041768f
C4853 VDPWR.n667 VGND 0.036489f
C4854 VDPWR.n668 VGND 0.041768f
C4855 VDPWR.n669 VGND 0.073918f
C4856 VDPWR.n670 VGND 0.046407f
C4857 VDPWR.n671 VGND 0.006601f
C4858 VDPWR.n672 VGND 0.503555f
C4859 VDPWR.n673 VGND 0.078633f
C4860 VDPWR.n674 VGND 0.078633f
C4861 VDPWR.n675 VGND 0.065925f
C4862 VDPWR.n676 VGND 0.107512f
C4863 VDPWR.n677 VGND 0.202734f
C4864 VDPWR.n678 VGND 0.149751f
C4865 VDPWR.n679 VGND 0.121863f
C4866 VDPWR.t185 VGND 0.66253f
C4867 VDPWR.n680 VGND 0.155747f
C4868 VDPWR.n681 VGND 0.371223f
C4869 VDPWR.n682 VGND 0.39542f
C4870 VDPWR.n683 VGND 0.041768f
C4871 VDPWR.n684 VGND 0.036489f
C4872 VDPWR.n685 VGND 0.041768f
C4873 VDPWR.n686 VGND 0.073918f
C4874 VDPWR.n687 VGND 0.046407f
C4875 VDPWR.n688 VGND 0.006601f
C4876 VDPWR.n689 VGND 0.503555f
C4877 VDPWR.n690 VGND 0.078633f
C4878 VDPWR.n691 VGND 0.078633f
C4879 VDPWR.n692 VGND 0.065925f
C4880 VDPWR.n693 VGND 0.107512f
C4881 VDPWR.n694 VGND 0.202734f
C4882 VDPWR.n695 VGND 0.149751f
C4883 VDPWR.n696 VGND 0.121863f
C4884 VDPWR.t118 VGND 0.66253f
C4885 VDPWR.n697 VGND 0.155747f
C4886 VDPWR.n698 VGND 0.371223f
C4887 VDPWR.n699 VGND 0.39542f
C4888 VDPWR.n700 VGND 0.041768f
C4889 VDPWR.n701 VGND 0.036489f
C4890 VDPWR.n702 VGND 0.041768f
C4891 VDPWR.n703 VGND 0.073918f
C4892 VDPWR.n704 VGND 0.046407f
C4893 VDPWR.n705 VGND 0.006601f
C4894 VDPWR.n706 VGND 0.503555f
C4895 VDPWR.n707 VGND 0.078633f
C4896 VDPWR.n708 VGND 0.078633f
C4897 VDPWR.n709 VGND 0.065925f
C4898 VDPWR.n710 VGND 0.107512f
C4899 VDPWR.n711 VGND 0.046716f
C4900 VDPWR.t107 VGND 0.050473f
C4901 VDPWR.n712 VGND 0.093119f
C4902 VDPWR.n713 VGND 0.041191f
C4903 VDPWR.n714 VGND 0.043552f
C4904 VDPWR.n715 VGND 0.021519f
C4905 VDPWR.n716 VGND 0.030925f
C4906 VDPWR.n717 VGND 0.051783f
C4907 VDPWR.t19 VGND 0.050473f
C4908 VDPWR.n718 VGND 0.043552f
C4909 VDPWR.t25 VGND 0.050473f
C4910 VDPWR.n719 VGND 0.093119f
C4911 VDPWR.n720 VGND 0.021519f
C4912 VDPWR.n721 VGND 0.043552f
C4913 VDPWR.n722 VGND 0.021519f
C4914 VDPWR.n723 VGND 0.030925f
C4915 VDPWR.n724 VGND 0.051783f
C4916 VDPWR.t27 VGND 0.050473f
C4917 VDPWR.n725 VGND 0.043552f
C4918 VDPWR.t22 VGND 0.050473f
C4919 VDPWR.n726 VGND 0.093119f
C4920 VDPWR.n727 VGND 0.021519f
C4921 VDPWR.n728 VGND 0.043552f
C4922 VDPWR.n729 VGND 0.021519f
C4923 VDPWR.n730 VGND 0.030925f
C4924 VDPWR.n731 VGND 0.051783f
C4925 VDPWR.t21 VGND 0.050473f
C4926 VDPWR.n732 VGND 0.043552f
C4927 VDPWR.t109 VGND 0.050473f
C4928 VDPWR.n733 VGND 0.093119f
C4929 VDPWR.n734 VGND 0.021519f
C4930 VDPWR.n735 VGND 0.043552f
C4931 VDPWR.n736 VGND 0.021519f
C4932 VDPWR.n737 VGND 0.030925f
C4933 VDPWR.n738 VGND 0.051783f
C4934 VDPWR.t111 VGND 0.050473f
C4935 VDPWR.n739 VGND 0.043552f
C4936 VDPWR.t24 VGND 0.050473f
C4937 VDPWR.n740 VGND 0.093119f
C4938 VDPWR.n741 VGND 0.021519f
C4939 VDPWR.n742 VGND 0.043552f
C4940 VDPWR.n743 VGND 0.021519f
C4941 VDPWR.n744 VGND 0.030925f
C4942 VDPWR.n745 VGND 0.051783f
C4943 VDPWR.t29 VGND 0.050473f
C4944 VDPWR.n746 VGND 0.043552f
C4945 VDPWR.t23 VGND 0.050473f
C4946 VDPWR.n747 VGND 0.093119f
C4947 VDPWR.n748 VGND 0.021519f
C4948 VDPWR.n749 VGND 0.043552f
C4949 VDPWR.n750 VGND 0.021519f
C4950 VDPWR.n751 VGND 0.030925f
C4951 VDPWR.n752 VGND 0.051783f
C4952 VDPWR.t28 VGND 0.050473f
C4953 VDPWR.n753 VGND 0.043552f
C4954 VDPWR.t20 VGND 0.050473f
C4955 VDPWR.n754 VGND 0.093119f
C4956 VDPWR.n755 VGND 0.021519f
C4957 VDPWR.n756 VGND 0.043552f
C4958 VDPWR.n757 VGND 0.021519f
C4959 VDPWR.n758 VGND 0.030925f
C4960 VDPWR.n759 VGND 0.051783f
C4961 VDPWR.t108 VGND 0.050473f
C4962 VDPWR.n760 VGND 0.043552f
C4963 VDPWR.t110 VGND 0.050473f
C4964 VDPWR.n761 VGND 0.093119f
C4965 VDPWR.n762 VGND 0.021519f
C4966 VDPWR.n763 VGND 0.043552f
C4967 VDPWR.n764 VGND 0.021519f
C4968 VDPWR.n765 VGND 0.030925f
C4969 VDPWR.n766 VGND 0.051783f
C4970 VDPWR.t26 VGND 0.050473f
C4971 VDPWR.n767 VGND 0.043552f
C4972 VDPWR.t596 VGND 0.050473f
C4973 VDPWR.n768 VGND 0.093119f
C4974 VDPWR.n769 VGND 0.021519f
C4975 VDPWR.n770 VGND 0.043552f
C4976 VDPWR.n771 VGND 0.021519f
C4977 VDPWR.n772 VGND 0.030925f
C4978 VDPWR.n773 VGND 0.051783f
C4979 VDPWR.t598 VGND 0.050473f
C4980 VDPWR.n774 VGND 0.043552f
C4981 VDPWR.t599 VGND 0.050473f
C4982 VDPWR.n775 VGND 0.093119f
C4983 VDPWR.n776 VGND 0.021519f
C4984 VDPWR.n777 VGND 0.043552f
C4985 VDPWR.n778 VGND 0.021519f
C4986 VDPWR.n779 VGND 0.030925f
C4987 VDPWR.n780 VGND 0.051783f
C4988 VDPWR.t597 VGND 0.050473f
C4989 VDPWR.n781 VGND 0.043552f
C4990 VDPWR.t193 VGND 0.050473f
C4991 VDPWR.n782 VGND 0.093119f
C4992 VDPWR.n783 VGND 0.021519f
C4993 VDPWR.n784 VGND 0.043552f
C4994 VDPWR.n785 VGND 0.021519f
C4995 VDPWR.n786 VGND 0.030925f
C4996 VDPWR.n787 VGND 0.051783f
C4997 VDPWR.t400 VGND 0.050473f
C4998 VDPWR.n788 VGND 0.043552f
C4999 VDPWR.t225 VGND 0.050473f
C5000 VDPWR.n789 VGND 0.093119f
C5001 VDPWR.n790 VGND 0.021519f
C5002 VDPWR.n791 VGND 0.043552f
C5003 VDPWR.n792 VGND 0.021519f
C5004 VDPWR.n793 VGND 0.030925f
C5005 VDPWR.n794 VGND 0.051783f
C5006 VDPWR.t290 VGND 0.050473f
C5007 VDPWR.n795 VGND 0.043552f
C5008 VDPWR.t164 VGND 0.050473f
C5009 VDPWR.n796 VGND 0.093119f
C5010 VDPWR.n797 VGND 0.021519f
C5011 VDPWR.n798 VGND 0.043552f
C5012 VDPWR.n799 VGND 0.021519f
C5013 VDPWR.n800 VGND 0.030925f
C5014 VDPWR.n801 VGND 0.051783f
C5015 VDPWR.t198 VGND 0.050473f
C5016 VDPWR.n802 VGND 0.043552f
C5017 VDPWR.t574 VGND 0.050473f
C5018 VDPWR.n803 VGND 0.093119f
C5019 VDPWR.n804 VGND 0.021519f
C5020 VDPWR.n805 VGND 0.043552f
C5021 VDPWR.n806 VGND 0.041191f
C5022 VDPWR.t18 VGND 4.75727f
C5023 VDPWR.n807 VGND 0.030825f
C5024 VDPWR.n808 VGND 0.030925f
C5025 VDPWR.n809 VGND 0.02766f
C5026 VDPWR.n810 VGND 0.030925f
C5027 VDPWR.n811 VGND 0.02766f
C5028 VDPWR.n812 VGND 0.030925f
C5029 VDPWR.n813 VGND 0.02766f
C5030 VDPWR.n814 VGND 0.030925f
C5031 VDPWR.n815 VGND 0.02766f
C5032 VDPWR.n816 VGND 0.030925f
C5033 VDPWR.n817 VGND 0.02766f
C5034 VDPWR.n818 VGND 0.030925f
C5035 VDPWR.n819 VGND 0.02766f
C5036 VDPWR.n820 VGND 0.030925f
C5037 VDPWR.n821 VGND 0.02766f
C5038 VDPWR.n822 VGND 0.030925f
C5039 VDPWR.n823 VGND 0.02766f
C5040 VDPWR.n824 VGND 0.030925f
C5041 VDPWR.n825 VGND 0.02766f
C5042 VDPWR.n826 VGND 0.030925f
C5043 VDPWR.n827 VGND 0.02766f
C5044 VDPWR.n828 VGND 0.030925f
C5045 VDPWR.n829 VGND 0.02766f
C5046 VDPWR.n830 VGND 0.030925f
C5047 VDPWR.n831 VGND 0.02766f
C5048 VDPWR.n832 VGND 0.030925f
C5049 VDPWR.n833 VGND 0.02766f
C5050 VDPWR.n834 VGND 0.030925f
C5051 VDPWR.n835 VGND 0.02766f
C5052 VDPWR.n836 VGND 0.030925f
C5053 VDPWR.n837 VGND 0.02766f
C5054 VDPWR.n838 VGND 0.030925f
C5055 VDPWR.n839 VGND 0.02766f
C5056 VDPWR.n840 VGND 0.030925f
C5057 VDPWR.n841 VGND 0.02766f
C5058 VDPWR.n842 VGND 0.030925f
C5059 VDPWR.n843 VGND 0.02766f
C5060 VDPWR.n844 VGND 0.030925f
C5061 VDPWR.n845 VGND 0.02766f
C5062 VDPWR.n846 VGND 0.030925f
C5063 VDPWR.n847 VGND 0.02766f
C5064 VDPWR.n848 VGND 0.030925f
C5065 VDPWR.n849 VGND 0.02766f
C5066 VDPWR.n850 VGND 0.030925f
C5067 VDPWR.n851 VGND 0.02766f
C5068 VDPWR.n852 VGND 0.030925f
C5069 VDPWR.n853 VGND 0.02766f
C5070 VDPWR.n854 VGND 0.030925f
C5071 VDPWR.n855 VGND 0.02766f
C5072 VDPWR.n856 VGND 0.030925f
C5073 VDPWR.n857 VGND 0.02766f
C5074 VDPWR.n858 VGND 0.030925f
C5075 VDPWR.n859 VGND 0.02766f
C5076 VDPWR.n860 VGND 3.52343f
C5077 VDPWR.n861 VGND 0.030925f
C5078 VDPWR.n862 VGND 0.02766f
C5079 VDPWR.n863 VGND 2.60759f
C5080 VDPWR.n864 VGND 0.030825f
C5081 VDPWR.n865 VGND 0.046716f
C5082 VDPWR.n866 VGND 0.051783f
C5083 VDPWR.t605 VGND 0.050473f
C5084 VDPWR.n867 VGND 0.045031f
C5085 VDPWR.n868 VGND 0.093119f
C5086 VDPWR.n869 VGND 0.014025f
C5087 VDPWR.n870 VGND 0.041191f
C5088 VDPWR.n871 VGND 0.030925f
C5089 VDPWR.n872 VGND 0.021519f
C5090 VDPWR.n873 VGND 0.014025f
C5091 VDPWR.n874 VGND 0.051783f
C5092 VDPWR.n875 VGND 0.093119f
C5093 VDPWR.n876 VGND 0.014025f
C5094 VDPWR.n877 VGND 0.021519f
C5095 VDPWR.n878 VGND 0.030925f
C5096 VDPWR.n879 VGND 0.021519f
C5097 VDPWR.n880 VGND 0.014025f
C5098 VDPWR.n881 VGND 0.051783f
C5099 VDPWR.n882 VGND 0.093119f
C5100 VDPWR.n883 VGND 0.014025f
C5101 VDPWR.n884 VGND 0.021519f
C5102 VDPWR.n885 VGND 0.030925f
C5103 VDPWR.n886 VGND 0.021519f
C5104 VDPWR.n887 VGND 0.014025f
C5105 VDPWR.n888 VGND 0.051783f
C5106 VDPWR.n889 VGND 0.093119f
C5107 VDPWR.n890 VGND 0.014025f
C5108 VDPWR.n891 VGND 0.021519f
C5109 VDPWR.n892 VGND 0.030925f
C5110 VDPWR.n893 VGND 0.021519f
C5111 VDPWR.n894 VGND 0.014025f
C5112 VDPWR.n895 VGND 0.051783f
C5113 VDPWR.n896 VGND 0.093119f
C5114 VDPWR.n897 VGND 0.014025f
C5115 VDPWR.n898 VGND 0.021519f
C5116 VDPWR.n899 VGND 0.030925f
C5117 VDPWR.n900 VGND 0.021519f
C5118 VDPWR.n901 VGND 0.014025f
C5119 VDPWR.n902 VGND 0.051783f
C5120 VDPWR.n903 VGND 0.093119f
C5121 VDPWR.n904 VGND 0.014025f
C5122 VDPWR.n905 VGND 0.021519f
C5123 VDPWR.n906 VGND 0.030925f
C5124 VDPWR.n907 VGND 0.021519f
C5125 VDPWR.n908 VGND 0.014025f
C5126 VDPWR.n909 VGND 0.051783f
C5127 VDPWR.n910 VGND 0.093119f
C5128 VDPWR.n911 VGND 0.014025f
C5129 VDPWR.n912 VGND 0.021519f
C5130 VDPWR.n913 VGND 0.030925f
C5131 VDPWR.n914 VGND 0.021519f
C5132 VDPWR.n915 VGND 0.014025f
C5133 VDPWR.n916 VGND 0.051783f
C5134 VDPWR.n917 VGND 0.093119f
C5135 VDPWR.n918 VGND 0.014025f
C5136 VDPWR.n919 VGND 0.021519f
C5137 VDPWR.n920 VGND 0.030925f
C5138 VDPWR.n921 VGND 0.021519f
C5139 VDPWR.n922 VGND 0.014025f
C5140 VDPWR.n923 VGND 0.051783f
C5141 VDPWR.n924 VGND 0.093119f
C5142 VDPWR.n925 VGND 0.014025f
C5143 VDPWR.n926 VGND 0.021519f
C5144 VDPWR.n927 VGND 0.030925f
C5145 VDPWR.n928 VGND 0.021519f
C5146 VDPWR.n929 VGND 0.014025f
C5147 VDPWR.n930 VGND 0.051783f
C5148 VDPWR.n931 VGND 0.093119f
C5149 VDPWR.n932 VGND 0.014025f
C5150 VDPWR.n933 VGND 0.021519f
C5151 VDPWR.n934 VGND 0.030925f
C5152 VDPWR.n935 VGND 0.021519f
C5153 VDPWR.n936 VGND 0.014025f
C5154 VDPWR.n937 VGND 0.051783f
C5155 VDPWR.n938 VGND 0.093119f
C5156 VDPWR.n939 VGND 0.014025f
C5157 VDPWR.n940 VGND 0.021519f
C5158 VDPWR.n941 VGND 0.030925f
C5159 VDPWR.n942 VGND 0.021519f
C5160 VDPWR.n943 VGND 0.014025f
C5161 VDPWR.n944 VGND 0.051783f
C5162 VDPWR.n945 VGND 0.093119f
C5163 VDPWR.n946 VGND 0.014025f
C5164 VDPWR.n947 VGND 0.021519f
C5165 VDPWR.n948 VGND 0.030925f
C5166 VDPWR.n949 VGND 0.021519f
C5167 VDPWR.n950 VGND 0.014025f
C5168 VDPWR.n951 VGND 0.051783f
C5169 VDPWR.n952 VGND 0.093119f
C5170 VDPWR.n953 VGND 0.014025f
C5171 VDPWR.n954 VGND 0.021519f
C5172 VDPWR.n955 VGND 0.030925f
C5173 VDPWR.n956 VGND 0.021519f
C5174 VDPWR.n957 VGND 0.014025f
C5175 VDPWR.n958 VGND 0.051783f
C5176 VDPWR.n959 VGND 0.093119f
C5177 VDPWR.n960 VGND 0.014025f
C5178 VDPWR.n961 VGND 0.021519f
C5179 VDPWR.n962 VGND 0.030925f
C5180 VDPWR.n963 VGND 0.041191f
C5181 VDPWR.n964 VGND 0.014025f
C5182 VDPWR.n965 VGND 0.09831f
C5183 VDPWR.n966 VGND 0.069174f
C5184 VDPWR.t318 VGND 0.01345f
C5185 VDPWR.t395 VGND 0.01345f
C5186 VDPWR.n967 VGND 0.028501f
C5187 VDPWR.t614 VGND 0.050702f
C5188 VDPWR.n968 VGND 0.049137f
C5189 VDPWR.t131 VGND 0.050702f
C5190 VDPWR.n969 VGND 0.116724f
C5191 VDPWR.n970 VGND 0.069174f
C5192 VDPWR.t513 VGND 0.01345f
C5193 VDPWR.t573 VGND 0.01345f
C5194 VDPWR.n971 VGND 0.028501f
C5195 VDPWR.t530 VGND 0.050702f
C5196 VDPWR.n972 VGND 0.049137f
C5197 VDPWR.t295 VGND 0.050702f
C5198 VDPWR.n973 VGND 0.116724f
C5199 VDPWR.n974 VGND 0.069174f
C5200 VDPWR.t537 VGND 0.01345f
C5201 VDPWR.t338 VGND 0.01345f
C5202 VDPWR.n975 VGND 0.028501f
C5203 VDPWR.t135 VGND 0.050702f
C5204 VDPWR.n976 VGND 0.049137f
C5205 VDPWR.t325 VGND 0.050702f
C5206 VDPWR.n977 VGND 0.116724f
C5207 VDPWR.n978 VGND 0.069174f
C5208 VDPWR.t539 VGND 0.01345f
C5209 VDPWR.t69 VGND 0.01345f
C5210 VDPWR.n979 VGND 0.028501f
C5211 VDPWR.t241 VGND 0.050702f
C5212 VDPWR.n980 VGND 0.049137f
C5213 VDPWR.t211 VGND 0.050702f
C5214 VDPWR.n981 VGND 0.116724f
C5215 VDPWR.n982 VGND 0.069174f
C5216 VDPWR.t63 VGND 0.01345f
C5217 VDPWR.t565 VGND 0.01345f
C5218 VDPWR.n983 VGND 0.028501f
C5219 VDPWR.t567 VGND 0.050702f
C5220 VDPWR.n984 VGND 0.049137f
C5221 VDPWR.t589 VGND 0.050702f
C5222 VDPWR.n985 VGND 0.116724f
C5223 VDPWR.n986 VGND 0.069174f
C5224 VDPWR.t347 VGND 0.01345f
C5225 VDPWR.t228 VGND 0.01345f
C5226 VDPWR.n987 VGND 0.028501f
C5227 VDPWR.t389 VGND 0.050702f
C5228 VDPWR.n988 VGND 0.049137f
C5229 VDPWR.t483 VGND 0.050702f
C5230 VDPWR.n989 VGND 0.116724f
C5231 VDPWR.n990 VGND 0.069174f
C5232 VDPWR.t620 VGND 0.01345f
C5233 VDPWR.t38 VGND 0.01345f
C5234 VDPWR.n991 VGND 0.028501f
C5235 VDPWR.t618 VGND 0.050702f
C5236 VDPWR.n992 VGND 0.049137f
C5237 VDPWR.t385 VGND 0.050702f
C5238 VDPWR.n993 VGND 0.116724f
C5239 VDPWR.n994 VGND 0.069174f
C5240 VDPWR.t102 VGND 0.01345f
C5241 VDPWR.t582 VGND 0.01345f
C5242 VDPWR.n995 VGND 0.028501f
C5243 VDPWR.t58 VGND 0.050702f
C5244 VDPWR.n996 VGND 0.049137f
C5245 VDPWR.t273 VGND 0.050702f
C5246 VDPWR.n997 VGND 0.116724f
C5247 VDPWR.t106 VGND 0.01345f
C5248 VDPWR.t213 VGND 0.01345f
C5249 VDPWR.n998 VGND 0.028501f
C5250 VDPWR.n999 VGND 0.24424f
C5251 VDPWR.n1000 VGND 0.082251f
C5252 VDPWR.n1001 VGND 0.265689f
C5253 VDPWR.n1002 VGND 0.100518f
C5254 VDPWR.t105 VGND 0.207052f
C5255 VDPWR.t212 VGND 0.130601f
C5256 VDPWR.t600 VGND 0.130601f
C5257 VDPWR.t272 VGND 0.171413f
C5258 VDPWR.n1003 VGND 0.263216f
C5259 VDPWR.t581 VGND 0.203489f
C5260 VDPWR.t101 VGND 0.130601f
C5261 VDPWR.t85 VGND 0.130601f
C5262 VDPWR.t57 VGND 0.172898f
C5263 VDPWR.n1004 VGND 0.029636f
C5264 VDPWR.n1005 VGND 0.109081f
C5265 VDPWR.n1006 VGND 0.107597f
C5266 VDPWR.n1007 VGND 0.088629f
C5267 VDPWR.n1008 VGND 0.100518f
C5268 VDPWR.n1009 VGND 0.088629f
C5269 VDPWR.n1010 VGND 0.007963f
C5270 VDPWR.n1011 VGND 0.044273f
C5271 VDPWR.n1012 VGND 0.116882f
C5272 VDPWR.n1013 VGND 0.119122f
C5273 VDPWR.n1014 VGND 0.058307f
C5274 VDPWR.t235 VGND 0.01345f
C5275 VDPWR.t97 VGND 0.01345f
C5276 VDPWR.n1015 VGND 0.028501f
C5277 VDPWR.n1016 VGND 0.119595f
C5278 VDPWR.n1017 VGND 0.094575f
C5279 VDPWR.n1018 VGND 0.069274f
C5280 VDPWR.n1019 VGND 0.265689f
C5281 VDPWR.n1020 VGND 0.100518f
C5282 VDPWR.t234 VGND 0.207052f
C5283 VDPWR.t96 VGND 0.130601f
C5284 VDPWR.t397 VGND 0.130601f
C5285 VDPWR.t384 VGND 0.171413f
C5286 VDPWR.n1021 VGND 0.263216f
C5287 VDPWR.t37 VGND 0.203489f
C5288 VDPWR.t619 VGND 0.130601f
C5289 VDPWR.t197 VGND 0.130601f
C5290 VDPWR.t617 VGND 0.172898f
C5291 VDPWR.n1022 VGND 0.029636f
C5292 VDPWR.n1023 VGND 0.109081f
C5293 VDPWR.n1024 VGND 0.107597f
C5294 VDPWR.n1025 VGND 0.088629f
C5295 VDPWR.n1026 VGND 0.100518f
C5296 VDPWR.n1027 VGND 0.088629f
C5297 VDPWR.n1028 VGND 0.007963f
C5298 VDPWR.n1029 VGND 0.044273f
C5299 VDPWR.n1030 VGND 0.116882f
C5300 VDPWR.n1031 VGND 0.119122f
C5301 VDPWR.n1032 VGND 0.058307f
C5302 VDPWR.t192 VGND 0.01345f
C5303 VDPWR.t230 VGND 0.01345f
C5304 VDPWR.n1033 VGND 0.028501f
C5305 VDPWR.n1034 VGND 0.119595f
C5306 VDPWR.n1035 VGND 0.094575f
C5307 VDPWR.n1036 VGND 0.069274f
C5308 VDPWR.n1037 VGND 0.265689f
C5309 VDPWR.n1038 VGND 0.100518f
C5310 VDPWR.t191 VGND 0.207052f
C5311 VDPWR.t229 VGND 0.130601f
C5312 VDPWR.t82 VGND 0.130601f
C5313 VDPWR.t482 VGND 0.171413f
C5314 VDPWR.n1039 VGND 0.263216f
C5315 VDPWR.t227 VGND 0.203489f
C5316 VDPWR.t346 VGND 0.130601f
C5317 VDPWR.t171 VGND 0.130601f
C5318 VDPWR.t388 VGND 0.172898f
C5319 VDPWR.n1040 VGND 0.029636f
C5320 VDPWR.n1041 VGND 0.109081f
C5321 VDPWR.n1042 VGND 0.107597f
C5322 VDPWR.n1043 VGND 0.088629f
C5323 VDPWR.n1044 VGND 0.100518f
C5324 VDPWR.n1045 VGND 0.088629f
C5325 VDPWR.n1046 VGND 0.007963f
C5326 VDPWR.n1047 VGND 0.044273f
C5327 VDPWR.n1048 VGND 0.116882f
C5328 VDPWR.n1049 VGND 0.119122f
C5329 VDPWR.n1050 VGND 0.058307f
C5330 VDPWR.t585 VGND 0.01345f
C5331 VDPWR.t563 VGND 0.01345f
C5332 VDPWR.n1051 VGND 0.028501f
C5333 VDPWR.n1052 VGND 0.119595f
C5334 VDPWR.n1053 VGND 0.094575f
C5335 VDPWR.n1054 VGND 0.069274f
C5336 VDPWR.n1055 VGND 0.265689f
C5337 VDPWR.n1056 VGND 0.100518f
C5338 VDPWR.t584 VGND 0.207052f
C5339 VDPWR.t562 VGND 0.130601f
C5340 VDPWR.t476 VGND 0.130601f
C5341 VDPWR.t588 VGND 0.171413f
C5342 VDPWR.n1057 VGND 0.263216f
C5343 VDPWR.t564 VGND 0.203489f
C5344 VDPWR.t62 VGND 0.130601f
C5345 VDPWR.t194 VGND 0.130601f
C5346 VDPWR.t566 VGND 0.172898f
C5347 VDPWR.n1058 VGND 0.029636f
C5348 VDPWR.n1059 VGND 0.109081f
C5349 VDPWR.n1060 VGND 0.107597f
C5350 VDPWR.n1061 VGND 0.088629f
C5351 VDPWR.n1062 VGND 0.100518f
C5352 VDPWR.n1063 VGND 0.088629f
C5353 VDPWR.n1064 VGND 0.007963f
C5354 VDPWR.n1065 VGND 0.044273f
C5355 VDPWR.n1066 VGND 0.116882f
C5356 VDPWR.n1067 VGND 0.119122f
C5357 VDPWR.n1068 VGND 0.058307f
C5358 VDPWR.t155 VGND 0.01345f
C5359 VDPWR.t201 VGND 0.01345f
C5360 VDPWR.n1069 VGND 0.028501f
C5361 VDPWR.n1070 VGND 0.119595f
C5362 VDPWR.n1071 VGND 0.094575f
C5363 VDPWR.n1072 VGND 0.069274f
C5364 VDPWR.n1073 VGND 0.265689f
C5365 VDPWR.n1074 VGND 0.100518f
C5366 VDPWR.t154 VGND 0.207052f
C5367 VDPWR.t200 VGND 0.130601f
C5368 VDPWR.t173 VGND 0.130601f
C5369 VDPWR.t210 VGND 0.171413f
C5370 VDPWR.n1075 VGND 0.263216f
C5371 VDPWR.t68 VGND 0.203489f
C5372 VDPWR.t538 VGND 0.130601f
C5373 VDPWR.t32 VGND 0.130601f
C5374 VDPWR.t240 VGND 0.172898f
C5375 VDPWR.n1076 VGND 0.029636f
C5376 VDPWR.n1077 VGND 0.109081f
C5377 VDPWR.n1078 VGND 0.107597f
C5378 VDPWR.n1079 VGND 0.088629f
C5379 VDPWR.n1080 VGND 0.100518f
C5380 VDPWR.n1081 VGND 0.088629f
C5381 VDPWR.n1082 VGND 0.007963f
C5382 VDPWR.n1083 VGND 0.044273f
C5383 VDPWR.n1084 VGND 0.116882f
C5384 VDPWR.n1085 VGND 0.119122f
C5385 VDPWR.n1086 VGND 0.058307f
C5386 VDPWR.t402 VGND 0.01345f
C5387 VDPWR.t336 VGND 0.01345f
C5388 VDPWR.n1087 VGND 0.028501f
C5389 VDPWR.n1088 VGND 0.119595f
C5390 VDPWR.n1089 VGND 0.094575f
C5391 VDPWR.n1090 VGND 0.069274f
C5392 VDPWR.n1091 VGND 0.265689f
C5393 VDPWR.n1092 VGND 0.100518f
C5394 VDPWR.t401 VGND 0.207052f
C5395 VDPWR.t335 VGND 0.130601f
C5396 VDPWR.t267 VGND 0.130601f
C5397 VDPWR.t324 VGND 0.171413f
C5398 VDPWR.n1093 VGND 0.263216f
C5399 VDPWR.t337 VGND 0.203489f
C5400 VDPWR.t536 VGND 0.130601f
C5401 VDPWR.t136 VGND 0.130601f
C5402 VDPWR.t134 VGND 0.172898f
C5403 VDPWR.n1094 VGND 0.029636f
C5404 VDPWR.n1095 VGND 0.109081f
C5405 VDPWR.n1096 VGND 0.107597f
C5406 VDPWR.n1097 VGND 0.088629f
C5407 VDPWR.n1098 VGND 0.100518f
C5408 VDPWR.n1099 VGND 0.088629f
C5409 VDPWR.n1100 VGND 0.007963f
C5410 VDPWR.n1101 VGND 0.044273f
C5411 VDPWR.n1102 VGND 0.116882f
C5412 VDPWR.n1103 VGND 0.119122f
C5413 VDPWR.n1104 VGND 0.058307f
C5414 VDPWR.t511 VGND 0.01345f
C5415 VDPWR.t345 VGND 0.01345f
C5416 VDPWR.n1105 VGND 0.028501f
C5417 VDPWR.n1106 VGND 0.119595f
C5418 VDPWR.n1107 VGND 0.094575f
C5419 VDPWR.n1108 VGND 0.069274f
C5420 VDPWR.n1109 VGND 0.265689f
C5421 VDPWR.n1110 VGND 0.100518f
C5422 VDPWR.t510 VGND 0.207052f
C5423 VDPWR.t344 VGND 0.130601f
C5424 VDPWR.t264 VGND 0.130601f
C5425 VDPWR.t294 VGND 0.171413f
C5426 VDPWR.n1111 VGND 0.263216f
C5427 VDPWR.t572 VGND 0.203489f
C5428 VDPWR.t512 VGND 0.130601f
C5429 VDPWR.t195 VGND 0.130601f
C5430 VDPWR.t529 VGND 0.172898f
C5431 VDPWR.n1112 VGND 0.029636f
C5432 VDPWR.n1113 VGND 0.109081f
C5433 VDPWR.n1114 VGND 0.107597f
C5434 VDPWR.n1115 VGND 0.088629f
C5435 VDPWR.n1116 VGND 0.100518f
C5436 VDPWR.n1117 VGND 0.088629f
C5437 VDPWR.n1118 VGND 0.007963f
C5438 VDPWR.n1119 VGND 0.044273f
C5439 VDPWR.n1120 VGND 0.116882f
C5440 VDPWR.n1121 VGND 0.119122f
C5441 VDPWR.n1122 VGND 0.058307f
C5442 VDPWR.t41 VGND 0.01345f
C5443 VDPWR.t117 VGND 0.01345f
C5444 VDPWR.n1123 VGND 0.028501f
C5445 VDPWR.n1124 VGND 0.119595f
C5446 VDPWR.n1125 VGND 0.094575f
C5447 VDPWR.n1126 VGND 0.069274f
C5448 VDPWR.n1127 VGND 0.265689f
C5449 VDPWR.n1128 VGND 0.100518f
C5450 VDPWR.t40 VGND 0.207052f
C5451 VDPWR.t116 VGND 0.130601f
C5452 VDPWR.t196 VGND 0.130601f
C5453 VDPWR.t130 VGND 0.171413f
C5454 VDPWR.n1129 VGND 0.263216f
C5455 VDPWR.t394 VGND 0.203489f
C5456 VDPWR.t317 VGND 0.130601f
C5457 VDPWR.t15 VGND 0.130601f
C5458 VDPWR.t613 VGND 0.172898f
C5459 VDPWR.n1130 VGND 0.029636f
C5460 VDPWR.n1131 VGND 0.109081f
C5461 VDPWR.n1132 VGND 0.107597f
C5462 VDPWR.n1133 VGND 0.088629f
C5463 VDPWR.n1134 VGND 0.100518f
C5464 VDPWR.n1135 VGND 0.088629f
C5465 VDPWR.n1136 VGND 0.007963f
C5466 VDPWR.n1137 VGND 0.044273f
C5467 VDPWR.n1138 VGND 0.116882f
C5468 VDPWR.n1139 VGND 0.119122f
C5469 VDPWR.n1140 VGND 0.058307f
C5470 VDPWR.n1141 VGND 0.544127f
C5471 VDPWR.n1142 VGND 0.318893f
C5472 VDPWR.n1143 VGND 0.077975f
C5473 VDPWR.t224 VGND 0.01345f
C5474 VDPWR.t133 VGND 0.01345f
C5475 VDPWR.n1144 VGND 0.028749f
C5476 VDPWR.t161 VGND 0.01345f
C5477 VDPWR.t602 VGND 0.01345f
C5478 VDPWR.n1145 VGND 0.028749f
C5479 VDPWR.t595 VGND 0.01345f
C5480 VDPWR.t50 VGND 0.01345f
C5481 VDPWR.n1146 VGND 0.028749f
C5482 VDPWR.n1147 VGND 0.116303f
C5483 VDPWR.n1148 VGND 0.077975f
C5484 VDPWR.t490 VGND 0.01345f
C5485 VDPWR.t383 VGND 0.01345f
C5486 VDPWR.n1149 VGND 0.028749f
C5487 VDPWR.t232 VGND 0.01345f
C5488 VDPWR.t492 VGND 0.01345f
C5489 VDPWR.n1150 VGND 0.028749f
C5490 VDPWR.t127 VGND 0.01345f
C5491 VDPWR.t54 VGND 0.01345f
C5492 VDPWR.n1151 VGND 0.028749f
C5493 VDPWR.n1152 VGND 0.116303f
C5494 VDPWR.n1153 VGND 0.077975f
C5495 VDPWR.t13 VGND 0.01345f
C5496 VDPWR.t7 VGND 0.01345f
C5497 VDPWR.n1154 VGND 0.028749f
C5498 VDPWR.t5 VGND 0.01345f
C5499 VDPWR.t239 VGND 0.01345f
C5500 VDPWR.n1155 VGND 0.028749f
C5501 VDPWR.t372 VGND 0.01345f
C5502 VDPWR.t370 VGND 0.01345f
C5503 VDPWR.n1156 VGND 0.028749f
C5504 VDPWR.n1157 VGND 0.116303f
C5505 VDPWR.n1158 VGND 0.077975f
C5506 VDPWR.t378 VGND 0.01345f
C5507 VDPWR.t360 VGND 0.01345f
C5508 VDPWR.n1159 VGND 0.028749f
C5509 VDPWR.t329 VGND 0.01345f
C5510 VDPWR.t362 VGND 0.01345f
C5511 VDPWR.n1160 VGND 0.028749f
C5512 VDPWR.t456 VGND 0.01345f
C5513 VDPWR.t458 VGND 0.01345f
C5514 VDPWR.n1161 VGND 0.028749f
C5515 VDPWR.n1162 VGND 0.116303f
C5516 VDPWR.n1163 VGND 0.077975f
C5517 VDPWR.t247 VGND 0.01345f
C5518 VDPWR.t168 VGND 0.01345f
C5519 VDPWR.n1164 VGND 0.028749f
C5520 VDPWR.t87 VGND 0.01345f
C5521 VDPWR.t499 VGND 0.01345f
C5522 VDPWR.n1165 VGND 0.028749f
C5523 VDPWR.t282 VGND 0.01345f
C5524 VDPWR.t280 VGND 0.01345f
C5525 VDPWR.n1166 VGND 0.028749f
C5526 VDPWR.n1167 VGND 0.116303f
C5527 VDPWR.n1168 VGND 0.077975f
C5528 VDPWR.t391 VGND 0.01345f
C5529 VDPWR.t163 VGND 0.01345f
C5530 VDPWR.n1169 VGND 0.028749f
C5531 VDPWR.t604 VGND 0.01345f
C5532 VDPWR.t60 VGND 0.01345f
C5533 VDPWR.n1170 VGND 0.028749f
C5534 VDPWR.t93 VGND 0.01345f
C5535 VDPWR.t578 VGND 0.01345f
C5536 VDPWR.n1171 VGND 0.028749f
C5537 VDPWR.n1172 VGND 0.116303f
C5538 VDPWR.n1173 VGND 0.077975f
C5539 VDPWR.t522 VGND 0.01345f
C5540 VDPWR.t31 VGND 0.01345f
C5541 VDPWR.n1174 VGND 0.028749f
C5542 VDPWR.t399 VGND 0.01345f
C5543 VDPWR.t524 VGND 0.01345f
C5544 VDPWR.n1175 VGND 0.028749f
C5545 VDPWR.t218 VGND 0.01345f
C5546 VDPWR.t207 VGND 0.01345f
C5547 VDPWR.n1176 VGND 0.028749f
C5548 VDPWR.n1177 VGND 0.116303f
C5549 VDPWR.n1178 VGND 0.077975f
C5550 VDPWR.t541 VGND 0.01345f
C5551 VDPWR.t587 VGND 0.01345f
C5552 VDPWR.n1179 VGND 0.028749f
C5553 VDPWR.t67 VGND 0.01345f
C5554 VDPWR.t65 VGND 0.01345f
C5555 VDPWR.n1180 VGND 0.028749f
C5556 VDPWR.t175 VGND 0.01345f
C5557 VDPWR.t190 VGND 0.01345f
C5558 VDPWR.n1181 VGND 0.028749f
C5559 VDPWR.n1182 VGND 0.116303f
C5560 VDPWR.n1183 VGND 0.078671f
C5561 VDPWR.t333 VGND 0.01345f
C5562 VDPWR.t331 VGND 0.01345f
C5563 VDPWR.n1184 VGND 0.028749f
C5564 VDPWR.t571 VGND 0.01345f
C5565 VDPWR.t269 VGND 0.01345f
C5566 VDPWR.n1185 VGND 0.028749f
C5567 VDPWR.t393 VGND 0.01345f
C5568 VDPWR.t350 VGND 0.01345f
C5569 VDPWR.n1186 VGND 0.028749f
C5570 VDPWR.n1187 VGND 0.116303f
C5571 VDPWR.n1188 VGND 0.094826f
C5572 VDPWR.n1189 VGND 0.090956f
C5573 VDPWR.n1190 VGND 0.052722f
C5574 VDPWR.t507 VGND 0.01345f
C5575 VDPWR.t466 VGND 0.01345f
C5576 VDPWR.n1191 VGND 0.028749f
C5577 VDPWR.n1192 VGND 0.167117f
C5578 VDPWR.n1193 VGND 0.085353f
C5579 VDPWR.n1194 VGND 0.230291f
C5580 VDPWR.t506 VGND 0.205794f
C5581 VDPWR.t465 VGND 0.138763f
C5582 VDPWR.t392 VGND 0.138763f
C5583 VDPWR.t349 VGND 0.184492f
C5584 VDPWR.n1195 VGND 0.068975f
C5585 VDPWR.n1196 VGND 0.118264f
C5586 VDPWR.n1197 VGND 0.156897f
C5587 VDPWR.t330 VGND 0.183704f
C5588 VDPWR.t332 VGND 0.138763f
C5589 VDPWR.t268 VGND 0.138763f
C5590 VDPWR.t570 VGND 0.181338f
C5591 VDPWR.n1198 VGND 0.11511f
C5592 VDPWR.n1199 VGND 0.078212f
C5593 VDPWR.n1200 VGND 0.078212f
C5594 VDPWR.n1201 VGND 0.028198f
C5595 VDPWR.n1202 VGND 0.115709f
C5596 VDPWR.n1203 VGND 0.115932f
C5597 VDPWR.n1204 VGND 0.136634f
C5598 VDPWR.t551 VGND 0.01345f
C5599 VDPWR.t177 VGND 0.01345f
C5600 VDPWR.n1205 VGND 0.028749f
C5601 VDPWR.n1206 VGND 0.115932f
C5602 VDPWR.n1207 VGND 0.136634f
C5603 VDPWR.n1208 VGND 0.077668f
C5604 VDPWR.n1209 VGND 0.169644f
C5605 VDPWR.n1210 VGND 0.229101f
C5606 VDPWR.t550 VGND 0.205794f
C5607 VDPWR.t176 VGND 0.138763f
C5608 VDPWR.t174 VGND 0.138763f
C5609 VDPWR.t189 VGND 0.184492f
C5610 VDPWR.n1211 VGND 0.052026f
C5611 VDPWR.n1212 VGND 0.156897f
C5612 VDPWR.t586 VGND 0.183704f
C5613 VDPWR.t540 VGND 0.138763f
C5614 VDPWR.t64 VGND 0.138763f
C5615 VDPWR.t66 VGND 0.181338f
C5616 VDPWR.n1213 VGND 0.11511f
C5617 VDPWR.n1214 VGND 0.18323f
C5618 VDPWR.n1215 VGND 0.007051f
C5619 VDPWR.n1216 VGND 0.173291f
C5620 VDPWR.n1217 VGND 0.028198f
C5621 VDPWR.n1218 VGND 0.115709f
C5622 VDPWR.n1219 VGND 0.115932f
C5623 VDPWR.n1220 VGND 0.136634f
C5624 VDPWR.t288 VGND 0.01345f
C5625 VDPWR.t297 VGND 0.01345f
C5626 VDPWR.n1221 VGND 0.028749f
C5627 VDPWR.n1222 VGND 0.115932f
C5628 VDPWR.n1223 VGND 0.136634f
C5629 VDPWR.n1224 VGND 0.077668f
C5630 VDPWR.n1225 VGND 0.169644f
C5631 VDPWR.n1226 VGND 0.229101f
C5632 VDPWR.t287 VGND 0.205794f
C5633 VDPWR.t296 VGND 0.138763f
C5634 VDPWR.t217 VGND 0.138763f
C5635 VDPWR.t206 VGND 0.184492f
C5636 VDPWR.n1227 VGND 0.052026f
C5637 VDPWR.n1228 VGND 0.156897f
C5638 VDPWR.t30 VGND 0.183704f
C5639 VDPWR.t521 VGND 0.138763f
C5640 VDPWR.t523 VGND 0.138763f
C5641 VDPWR.t398 VGND 0.181338f
C5642 VDPWR.n1229 VGND 0.11511f
C5643 VDPWR.n1230 VGND 0.18323f
C5644 VDPWR.n1231 VGND 0.007051f
C5645 VDPWR.n1232 VGND 0.173291f
C5646 VDPWR.n1233 VGND 0.028198f
C5647 VDPWR.n1234 VGND 0.115709f
C5648 VDPWR.n1235 VGND 0.115932f
C5649 VDPWR.n1236 VGND 0.136634f
C5650 VDPWR.t411 VGND 0.01345f
C5651 VDPWR.t48 VGND 0.01345f
C5652 VDPWR.n1237 VGND 0.028749f
C5653 VDPWR.n1238 VGND 0.115932f
C5654 VDPWR.n1239 VGND 0.136634f
C5655 VDPWR.n1240 VGND 0.077668f
C5656 VDPWR.n1241 VGND 0.169644f
C5657 VDPWR.n1242 VGND 0.229101f
C5658 VDPWR.t410 VGND 0.205794f
C5659 VDPWR.t47 VGND 0.138763f
C5660 VDPWR.t92 VGND 0.138763f
C5661 VDPWR.t577 VGND 0.184492f
C5662 VDPWR.n1243 VGND 0.052026f
C5663 VDPWR.n1244 VGND 0.156897f
C5664 VDPWR.t162 VGND 0.183704f
C5665 VDPWR.t390 VGND 0.138763f
C5666 VDPWR.t59 VGND 0.138763f
C5667 VDPWR.t603 VGND 0.181338f
C5668 VDPWR.n1245 VGND 0.11511f
C5669 VDPWR.n1246 VGND 0.18323f
C5670 VDPWR.n1247 VGND 0.007051f
C5671 VDPWR.n1248 VGND 0.173291f
C5672 VDPWR.n1249 VGND 0.028198f
C5673 VDPWR.n1250 VGND 0.115709f
C5674 VDPWR.n1251 VGND 0.115932f
C5675 VDPWR.n1252 VGND 0.136634f
C5676 VDPWR.t183 VGND 0.01345f
C5677 VDPWR.t481 VGND 0.01345f
C5678 VDPWR.n1253 VGND 0.028749f
C5679 VDPWR.n1254 VGND 0.115932f
C5680 VDPWR.n1255 VGND 0.136634f
C5681 VDPWR.n1256 VGND 0.077668f
C5682 VDPWR.n1257 VGND 0.169644f
C5683 VDPWR.n1258 VGND 0.229101f
C5684 VDPWR.t182 VGND 0.205794f
C5685 VDPWR.t480 VGND 0.138763f
C5686 VDPWR.t281 VGND 0.138763f
C5687 VDPWR.t279 VGND 0.184492f
C5688 VDPWR.n1259 VGND 0.052026f
C5689 VDPWR.n1260 VGND 0.156897f
C5690 VDPWR.t167 VGND 0.183704f
C5691 VDPWR.t246 VGND 0.138763f
C5692 VDPWR.t498 VGND 0.138763f
C5693 VDPWR.t86 VGND 0.181338f
C5694 VDPWR.n1261 VGND 0.11511f
C5695 VDPWR.n1262 VGND 0.18323f
C5696 VDPWR.n1263 VGND 0.007051f
C5697 VDPWR.n1264 VGND 0.173291f
C5698 VDPWR.n1265 VGND 0.028198f
C5699 VDPWR.n1266 VGND 0.115709f
C5700 VDPWR.n1267 VGND 0.115932f
C5701 VDPWR.n1268 VGND 0.136634f
C5702 VDPWR.t460 VGND 0.01345f
C5703 VDPWR.t454 VGND 0.01345f
C5704 VDPWR.n1269 VGND 0.028749f
C5705 VDPWR.n1270 VGND 0.115932f
C5706 VDPWR.n1271 VGND 0.136634f
C5707 VDPWR.n1272 VGND 0.077668f
C5708 VDPWR.n1273 VGND 0.169644f
C5709 VDPWR.n1274 VGND 0.229101f
C5710 VDPWR.t459 VGND 0.205794f
C5711 VDPWR.t453 VGND 0.138763f
C5712 VDPWR.t455 VGND 0.138763f
C5713 VDPWR.t457 VGND 0.184492f
C5714 VDPWR.n1275 VGND 0.052026f
C5715 VDPWR.n1276 VGND 0.156897f
C5716 VDPWR.t359 VGND 0.183704f
C5717 VDPWR.t377 VGND 0.138763f
C5718 VDPWR.t361 VGND 0.138763f
C5719 VDPWR.t328 VGND 0.181338f
C5720 VDPWR.n1277 VGND 0.11511f
C5721 VDPWR.n1278 VGND 0.18323f
C5722 VDPWR.n1279 VGND 0.007051f
C5723 VDPWR.n1280 VGND 0.173291f
C5724 VDPWR.n1281 VGND 0.028198f
C5725 VDPWR.n1282 VGND 0.115709f
C5726 VDPWR.n1283 VGND 0.115932f
C5727 VDPWR.n1284 VGND 0.136634f
C5728 VDPWR.t113 VGND 0.01345f
C5729 VDPWR.t409 VGND 0.01345f
C5730 VDPWR.n1285 VGND 0.028749f
C5731 VDPWR.n1286 VGND 0.115932f
C5732 VDPWR.n1287 VGND 0.136634f
C5733 VDPWR.n1288 VGND 0.077668f
C5734 VDPWR.n1289 VGND 0.169644f
C5735 VDPWR.n1290 VGND 0.229101f
C5736 VDPWR.t112 VGND 0.205794f
C5737 VDPWR.t408 VGND 0.138763f
C5738 VDPWR.t371 VGND 0.138763f
C5739 VDPWR.t369 VGND 0.184492f
C5740 VDPWR.n1291 VGND 0.052026f
C5741 VDPWR.n1292 VGND 0.156897f
C5742 VDPWR.t6 VGND 0.183704f
C5743 VDPWR.t12 VGND 0.138763f
C5744 VDPWR.t238 VGND 0.138763f
C5745 VDPWR.t4 VGND 0.181338f
C5746 VDPWR.n1293 VGND 0.11511f
C5747 VDPWR.n1294 VGND 0.18323f
C5748 VDPWR.n1295 VGND 0.007051f
C5749 VDPWR.n1296 VGND 0.173291f
C5750 VDPWR.n1297 VGND 0.028198f
C5751 VDPWR.n1298 VGND 0.115709f
C5752 VDPWR.n1299 VGND 0.115932f
C5753 VDPWR.n1300 VGND 0.136634f
C5754 VDPWR.t56 VGND 0.01345f
C5755 VDPWR.t505 VGND 0.01345f
C5756 VDPWR.n1301 VGND 0.028749f
C5757 VDPWR.n1302 VGND 0.115932f
C5758 VDPWR.n1303 VGND 0.136634f
C5759 VDPWR.n1304 VGND 0.077668f
C5760 VDPWR.n1305 VGND 0.169644f
C5761 VDPWR.n1306 VGND 0.229101f
C5762 VDPWR.t55 VGND 0.205794f
C5763 VDPWR.t504 VGND 0.138763f
C5764 VDPWR.t126 VGND 0.138763f
C5765 VDPWR.t53 VGND 0.184492f
C5766 VDPWR.n1307 VGND 0.052026f
C5767 VDPWR.n1308 VGND 0.156897f
C5768 VDPWR.t382 VGND 0.183704f
C5769 VDPWR.t489 VGND 0.138763f
C5770 VDPWR.t491 VGND 0.138763f
C5771 VDPWR.t231 VGND 0.181338f
C5772 VDPWR.n1309 VGND 0.11511f
C5773 VDPWR.n1310 VGND 0.18323f
C5774 VDPWR.n1311 VGND 0.007051f
C5775 VDPWR.n1312 VGND 0.173291f
C5776 VDPWR.n1313 VGND 0.028198f
C5777 VDPWR.n1314 VGND 0.115709f
C5778 VDPWR.n1315 VGND 0.115932f
C5779 VDPWR.n1316 VGND 0.136634f
C5780 VDPWR.t299 VGND 0.01345f
C5781 VDPWR.t263 VGND 0.01345f
C5782 VDPWR.n1317 VGND 0.028749f
C5783 VDPWR.n1318 VGND 0.115932f
C5784 VDPWR.n1319 VGND 0.136634f
C5785 VDPWR.n1320 VGND 0.077668f
C5786 VDPWR.n1321 VGND 0.169644f
C5787 VDPWR.n1322 VGND 0.229101f
C5788 VDPWR.t298 VGND 0.205794f
C5789 VDPWR.t262 VGND 0.138763f
C5790 VDPWR.t594 VGND 0.138763f
C5791 VDPWR.t49 VGND 0.184492f
C5792 VDPWR.n1323 VGND 0.052026f
C5793 VDPWR.n1324 VGND 0.156897f
C5794 VDPWR.t132 VGND 0.183704f
C5795 VDPWR.t223 VGND 0.138763f
C5796 VDPWR.t601 VGND 0.138763f
C5797 VDPWR.t160 VGND 0.181338f
C5798 VDPWR.n1325 VGND 0.11511f
C5799 VDPWR.n1326 VGND 0.18323f
C5800 VDPWR.n1327 VGND 0.007051f
C5801 VDPWR.n1328 VGND 0.173291f
C5802 VDPWR.n1329 VGND 0.028198f
C5803 VDPWR.n1330 VGND 0.115709f
C5804 VDPWR.n1331 VGND 0.115932f
C5805 VDPWR.n1332 VGND 0.09597f
C5806 VDPWR.n1333 VGND 0.228477f
C5807 VDPWR.n1334 VGND 6.55212f
C5808 VDPWR.n1335 VGND 0.077975f
C5809 VDPWR.t46 VGND 0.01345f
C5810 VDPWR.t404 VGND 0.01345f
C5811 VDPWR.n1336 VGND 0.028749f
C5812 VDPWR.t36 VGND 0.01345f
C5813 VDPWR.t44 VGND 0.01345f
C5814 VDPWR.n1337 VGND 0.028749f
C5815 VDPWR.t249 VGND 0.01345f
C5816 VDPWR.t251 VGND 0.01345f
C5817 VDPWR.n1338 VGND 0.028749f
C5818 VDPWR.n1339 VGND 0.116303f
C5819 VDPWR.n1340 VGND 0.077668f
C5820 VDPWR.n1341 VGND 0.169644f
C5821 VDPWR.t180 VGND 0.183704f
C5822 VDPWR.n1342 VGND 0.169951f
C5823 VDPWR.t253 VGND 0.01345f
C5824 VDPWR.t91 VGND 0.01345f
C5825 VDPWR.n1343 VGND 0.028749f
C5826 VDPWR.n1344 VGND 0.115932f
C5827 VDPWR.n1345 VGND 0.062281f
C5828 VDPWR.n1346 VGND 0.062281f
C5829 VDPWR.n1347 VGND 0.077668f
C5830 VDPWR.n1348 VGND 0.007051f
C5831 VDPWR.t501 VGND 0.01345f
C5832 VDPWR.t73 VGND 0.01345f
C5833 VDPWR.n1349 VGND 0.028749f
C5834 VDPWR.t129 VGND 0.01345f
C5835 VDPWR.t271 VGND 0.01345f
C5836 VDPWR.n1350 VGND 0.028749f
C5837 VDPWR.n1351 VGND 0.077668f
C5838 VDPWR.t220 VGND 0.01345f
C5839 VDPWR.t520 VGND 0.01345f
C5840 VDPWR.n1352 VGND 0.028749f
C5841 VDPWR.t495 VGND 0.01345f
C5842 VDPWR.t616 VGND 0.01345f
C5843 VDPWR.n1353 VGND 0.028749f
C5844 VDPWR.t374 VGND 0.01345f
C5845 VDPWR.t543 VGND 0.01345f
C5846 VDPWR.n1354 VGND 0.028749f
C5847 VDPWR.n1355 VGND 0.116303f
C5848 VDPWR.n1356 VGND 0.077668f
C5849 VDPWR.n1357 VGND 0.169951f
C5850 VDPWR.t471 VGND 0.183704f
C5851 VDPWR.n1358 VGND 0.169951f
C5852 VDPWR.t321 VGND 0.01345f
C5853 VDPWR.t140 VGND 0.01345f
C5854 VDPWR.n1359 VGND 0.028749f
C5855 VDPWR.n1360 VGND 0.115932f
C5856 VDPWR.n1361 VGND 0.062281f
C5857 VDPWR.n1362 VGND 0.062281f
C5858 VDPWR.n1363 VGND 0.077668f
C5859 VDPWR.n1364 VGND 0.007051f
C5860 VDPWR.t237 VGND 0.01345f
C5861 VDPWR.t209 VGND 0.01345f
C5862 VDPWR.n1365 VGND 0.028749f
C5863 VDPWR.t488 VGND 0.01345f
C5864 VDPWR.t464 VGND 0.01345f
C5865 VDPWR.n1366 VGND 0.028749f
C5866 VDPWR.n1367 VGND 0.077668f
C5867 VDPWR.t387 VGND 0.01345f
C5868 VDPWR.t144 VGND 0.01345f
C5869 VDPWR.n1368 VGND 0.028749f
C5870 VDPWR.t545 VGND 0.01345f
C5871 VDPWR.t323 VGND 0.01345f
C5872 VDPWR.n1369 VGND 0.028749f
C5873 VDPWR.t261 VGND 0.01345f
C5874 VDPWR.t561 VGND 0.01345f
C5875 VDPWR.n1370 VGND 0.028749f
C5876 VDPWR.n1371 VGND 0.116303f
C5877 VDPWR.n1372 VGND 0.077668f
C5878 VDPWR.n1373 VGND 0.169951f
C5879 VDPWR.t311 VGND 0.183704f
C5880 VDPWR.n1374 VGND 0.169951f
C5881 VDPWR.t559 VGND 0.01345f
C5882 VDPWR.t557 VGND 0.01345f
C5883 VDPWR.n1375 VGND 0.028749f
C5884 VDPWR.n1376 VGND 0.115932f
C5885 VDPWR.n1377 VGND 0.062281f
C5886 VDPWR.n1378 VGND 0.062281f
C5887 VDPWR.n1379 VGND 0.077668f
C5888 VDPWR.n1380 VGND 0.007051f
C5889 VDPWR.t591 VGND 0.01345f
C5890 VDPWR.t314 VGND 0.01345f
C5891 VDPWR.n1381 VGND 0.028749f
C5892 VDPWR.t316 VGND 0.01345f
C5893 VDPWR.t142 VGND 0.01345f
C5894 VDPWR.n1382 VGND 0.028749f
C5895 VDPWR.n1383 VGND 0.078671f
C5896 VDPWR.t9 VGND 0.01345f
C5897 VDPWR.t34 VGND 0.01345f
C5898 VDPWR.n1384 VGND 0.028749f
C5899 VDPWR.t147 VGND 0.01345f
C5900 VDPWR.t11 VGND 0.01345f
C5901 VDPWR.n1385 VGND 0.028749f
C5902 VDPWR.t376 VGND 0.01345f
C5903 VDPWR.t518 VGND 0.01345f
C5904 VDPWR.n1386 VGND 0.028749f
C5905 VDPWR.n1387 VGND 0.114596f
C5906 VDPWR.n1388 VGND 0.094826f
C5907 VDPWR.n1389 VGND 0.090956f
C5908 VDPWR.n1390 VGND 0.052722f
C5909 VDPWR.t159 VGND 0.01345f
C5910 VDPWR.t526 VGND 0.01345f
C5911 VDPWR.n1391 VGND 0.028905f
C5912 VDPWR.n1392 VGND 0.117409f
C5913 VDPWR.n1393 VGND 0.060979f
C5914 VDPWR.n1394 VGND 0.081124f
C5915 VDPWR.n1395 VGND 0.230291f
C5916 VDPWR.t158 VGND 0.205794f
C5917 VDPWR.t525 VGND 0.138763f
C5918 VDPWR.t375 VGND 0.138763f
C5919 VDPWR.t517 VGND 0.184492f
C5920 VDPWR.n1396 VGND 0.068975f
C5921 VDPWR.n1397 VGND 0.118264f
C5922 VDPWR.t496 VGND 0.138763f
C5923 VDPWR.t309 VGND 0.138763f
C5924 VDPWR.t307 VGND 0.181338f
C5925 VDPWR.n1398 VGND 0.11511f
C5926 VDPWR.n1399 VGND 0.18323f
C5927 VDPWR.t313 VGND 0.184492f
C5928 VDPWR.t590 VGND 0.138763f
C5929 VDPWR.t141 VGND 0.138763f
C5930 VDPWR.t315 VGND 0.183704f
C5931 VDPWR.n1400 VGND 0.051719f
C5932 VDPWR.n1401 VGND 0.20578f
C5933 VDPWR.n1402 VGND 0.156897f
C5934 VDPWR.t33 VGND 0.183704f
C5935 VDPWR.t8 VGND 0.138763f
C5936 VDPWR.t10 VGND 0.138763f
C5937 VDPWR.t146 VGND 0.181338f
C5938 VDPWR.n1403 VGND 0.11511f
C5939 VDPWR.n1404 VGND 0.078212f
C5940 VDPWR.n1405 VGND 0.078212f
C5941 VDPWR.n1406 VGND 0.028198f
C5942 VDPWR.n1407 VGND 0.115709f
C5943 VDPWR.n1408 VGND 0.115932f
C5944 VDPWR.n1409 VGND 0.062281f
C5945 VDPWR.n1410 VGND 0.062281f
C5946 VDPWR.n1411 VGND 0.115932f
C5947 VDPWR.n1412 VGND 0.116303f
C5948 VDPWR.t308 VGND 0.01345f
C5949 VDPWR.t310 VGND 0.01345f
C5950 VDPWR.n1413 VGND 0.028749f
C5951 VDPWR.t497 VGND 0.01345f
C5952 VDPWR.t312 VGND 0.01345f
C5953 VDPWR.n1414 VGND 0.028749f
C5954 VDPWR.n1415 VGND 0.115932f
C5955 VDPWR.n1416 VGND 0.115709f
C5956 VDPWR.n1417 VGND 0.028198f
C5957 VDPWR.n1418 VGND 0.173599f
C5958 VDPWR.n1419 VGND 0.077668f
C5959 VDPWR.n1420 VGND 0.051719f
C5960 VDPWR.n1421 VGND 0.156897f
C5961 VDPWR.n1422 VGND 0.051719f
C5962 VDPWR.n1423 VGND 0.20578f
C5963 VDPWR.t558 VGND 0.183704f
C5964 VDPWR.t556 VGND 0.138763f
C5965 VDPWR.t260 VGND 0.138763f
C5966 VDPWR.t560 VGND 0.184492f
C5967 VDPWR.t365 VGND 0.138763f
C5968 VDPWR.t367 VGND 0.138763f
C5969 VDPWR.t363 VGND 0.181338f
C5970 VDPWR.n1424 VGND 0.11511f
C5971 VDPWR.n1425 VGND 0.18323f
C5972 VDPWR.t208 VGND 0.184492f
C5973 VDPWR.t236 VGND 0.138763f
C5974 VDPWR.t463 VGND 0.138763f
C5975 VDPWR.t487 VGND 0.183704f
C5976 VDPWR.n1426 VGND 0.051719f
C5977 VDPWR.n1427 VGND 0.20578f
C5978 VDPWR.n1428 VGND 0.051719f
C5979 VDPWR.n1429 VGND 0.156897f
C5980 VDPWR.t143 VGND 0.183704f
C5981 VDPWR.t386 VGND 0.138763f
C5982 VDPWR.t322 VGND 0.138763f
C5983 VDPWR.t544 VGND 0.181338f
C5984 VDPWR.n1430 VGND 0.11511f
C5985 VDPWR.n1431 VGND 0.18323f
C5986 VDPWR.n1432 VGND 0.007051f
C5987 VDPWR.n1433 VGND 0.173599f
C5988 VDPWR.n1434 VGND 0.028198f
C5989 VDPWR.n1435 VGND 0.115709f
C5990 VDPWR.n1436 VGND 0.115932f
C5991 VDPWR.n1437 VGND 0.062281f
C5992 VDPWR.n1438 VGND 0.062281f
C5993 VDPWR.n1439 VGND 0.115932f
C5994 VDPWR.n1440 VGND 0.116303f
C5995 VDPWR.t364 VGND 0.01345f
C5996 VDPWR.t368 VGND 0.01345f
C5997 VDPWR.n1441 VGND 0.028749f
C5998 VDPWR.t366 VGND 0.01345f
C5999 VDPWR.t472 VGND 0.01345f
C6000 VDPWR.n1442 VGND 0.028749f
C6001 VDPWR.n1443 VGND 0.115932f
C6002 VDPWR.n1444 VGND 0.115709f
C6003 VDPWR.n1445 VGND 0.028198f
C6004 VDPWR.n1446 VGND 0.173599f
C6005 VDPWR.n1447 VGND 0.077668f
C6006 VDPWR.n1448 VGND 0.051719f
C6007 VDPWR.n1449 VGND 0.156897f
C6008 VDPWR.n1450 VGND 0.051719f
C6009 VDPWR.n1451 VGND 0.20578f
C6010 VDPWR.t320 VGND 0.183704f
C6011 VDPWR.t139 VGND 0.138763f
C6012 VDPWR.t373 VGND 0.138763f
C6013 VDPWR.t542 VGND 0.184492f
C6014 VDPWR.t467 VGND 0.138763f
C6015 VDPWR.t469 VGND 0.138763f
C6016 VDPWR.t178 VGND 0.181338f
C6017 VDPWR.n1452 VGND 0.11511f
C6018 VDPWR.n1453 VGND 0.18323f
C6019 VDPWR.t72 VGND 0.184492f
C6020 VDPWR.t500 VGND 0.138763f
C6021 VDPWR.t270 VGND 0.138763f
C6022 VDPWR.t128 VGND 0.183704f
C6023 VDPWR.n1454 VGND 0.051719f
C6024 VDPWR.n1455 VGND 0.20578f
C6025 VDPWR.n1456 VGND 0.051719f
C6026 VDPWR.n1457 VGND 0.156897f
C6027 VDPWR.t519 VGND 0.183704f
C6028 VDPWR.t219 VGND 0.138763f
C6029 VDPWR.t615 VGND 0.138763f
C6030 VDPWR.t494 VGND 0.181338f
C6031 VDPWR.n1458 VGND 0.11511f
C6032 VDPWR.n1459 VGND 0.18323f
C6033 VDPWR.n1460 VGND 0.007051f
C6034 VDPWR.n1461 VGND 0.173599f
C6035 VDPWR.n1462 VGND 0.028198f
C6036 VDPWR.n1463 VGND 0.115709f
C6037 VDPWR.n1464 VGND 0.115932f
C6038 VDPWR.n1465 VGND 0.062281f
C6039 VDPWR.n1466 VGND 0.062281f
C6040 VDPWR.n1467 VGND 0.115932f
C6041 VDPWR.n1468 VGND 0.116303f
C6042 VDPWR.t179 VGND 0.01345f
C6043 VDPWR.t470 VGND 0.01345f
C6044 VDPWR.n1469 VGND 0.028749f
C6045 VDPWR.t468 VGND 0.01345f
C6046 VDPWR.t181 VGND 0.01345f
C6047 VDPWR.n1470 VGND 0.028749f
C6048 VDPWR.n1471 VGND 0.115932f
C6049 VDPWR.n1472 VGND 0.115709f
C6050 VDPWR.n1473 VGND 0.028198f
C6051 VDPWR.n1474 VGND 0.173599f
C6052 VDPWR.n1475 VGND 0.077668f
C6053 VDPWR.n1476 VGND 0.051719f
C6054 VDPWR.n1477 VGND 0.156897f
C6055 VDPWR.n1478 VGND 0.051719f
C6056 VDPWR.n1479 VGND 0.20578f
C6057 VDPWR.t252 VGND 0.183704f
C6058 VDPWR.t90 VGND 0.138763f
C6059 VDPWR.t248 VGND 0.138763f
C6060 VDPWR.t250 VGND 0.184492f
C6061 VDPWR.n1480 VGND 0.052026f
C6062 VDPWR.n1481 VGND 0.156897f
C6063 VDPWR.t403 VGND 0.183704f
C6064 VDPWR.t45 VGND 0.138763f
C6065 VDPWR.t43 VGND 0.138763f
C6066 VDPWR.t35 VGND 0.181338f
C6067 VDPWR.n1482 VGND 0.11511f
C6068 VDPWR.n1483 VGND 0.18323f
C6069 VDPWR.n1484 VGND 0.007051f
C6070 VDPWR.n1485 VGND 0.173291f
C6071 VDPWR.n1486 VGND 0.028198f
C6072 VDPWR.n1487 VGND 0.115709f
C6073 VDPWR.n1488 VGND 0.115932f
C6074 VDPWR.n1489 VGND 0.058274f
C6075 VDPWR.n1490 VGND 0.046716f
C6076 VDPWR.t284 VGND 0.050473f
C6077 VDPWR.n1491 VGND 0.093119f
C6078 VDPWR.n1492 VGND 0.041191f
C6079 VDPWR.n1493 VGND 0.043552f
C6080 VDPWR.n1494 VGND 0.021519f
C6081 VDPWR.n1495 VGND 0.030925f
C6082 VDPWR.n1496 VGND 0.051783f
C6083 VDPWR.t172 VGND 0.050473f
C6084 VDPWR.n1497 VGND 0.043552f
C6085 VDPWR.t89 VGND 0.050473f
C6086 VDPWR.n1498 VGND 0.093119f
C6087 VDPWR.n1499 VGND 0.021519f
C6088 VDPWR.n1500 VGND 0.043552f
C6089 VDPWR.n1501 VGND 0.021519f
C6090 VDPWR.n1502 VGND 0.030925f
C6091 VDPWR.n1503 VGND 0.051783f
C6092 VDPWR.t302 VGND 0.050473f
C6093 VDPWR.n1504 VGND 0.043552f
C6094 VDPWR.t304 VGND 0.050473f
C6095 VDPWR.n1505 VGND 0.093119f
C6096 VDPWR.n1506 VGND 0.021519f
C6097 VDPWR.n1507 VGND 0.043552f
C6098 VDPWR.n1508 VGND 0.021519f
C6099 VDPWR.n1509 VGND 0.030925f
C6100 VDPWR.n1510 VGND 0.051783f
C6101 VDPWR.t301 VGND 0.050473f
C6102 VDPWR.n1511 VGND 0.010537f
C6103 VDPWR.n1512 VGND 0.030925f
C6104 VDPWR.t88 VGND 1.40382f
C6105 VDPWR.n1513 VGND 0.030825f
C6106 VDPWR.n1514 VGND 0.030925f
C6107 VDPWR.n1515 VGND 0.02766f
C6108 VDPWR.n1516 VGND 0.030925f
C6109 VDPWR.n1517 VGND 0.02766f
C6110 VDPWR.n1518 VGND 0.030925f
C6111 VDPWR.n1519 VGND 0.02766f
C6112 VDPWR.n1520 VGND 0.030925f
C6113 VDPWR.n1521 VGND 0.02766f
C6114 VDPWR.n1522 VGND 0.030925f
C6115 VDPWR.n1523 VGND 0.02766f
C6116 VDPWR.n1524 VGND 0.030825f
C6117 VDPWR.n1525 VGND 1.03973f
C6118 VDPWR.n1526 VGND 0.030925f
C6119 VDPWR.t303 VGND 0.050602f
C6120 VDPWR.n1527 VGND 0.094623f
C6121 VDPWR.n1528 VGND 0.051602f
C6122 VDPWR.n1529 VGND 0.021519f
C6123 VDPWR.n1530 VGND 0.021519f
C6124 VDPWR.n1531 VGND 0.041191f
C6125 VDPWR.n1532 VGND 0.048752f
C6126 VDPWR.n1533 VGND 0.044182f
C6127 VDPWR.t568 VGND 0.050602f
C6128 VDPWR.n1534 VGND 0.094623f
C6129 VDPWR.n1535 VGND 0.010537f
C6130 VDPWR.n1536 VGND 0.041191f
C6131 VDPWR.n1537 VGND 0.030925f
C6132 VDPWR.n1538 VGND 0.045588f
C6133 VDPWR.n1539 VGND 0.02766f
C6134 VDPWR.n1540 VGND 0.769474f
C6135 VDPWR.n1541 VGND 0.02766f
C6136 VDPWR.n1542 VGND 0.045588f
C6137 VDPWR.n1543 VGND 0.053309f
C6138 VDPWR.n1544 VGND 0.091339f
C6139 VDPWR.n1545 VGND 0.014025f
C6140 VDPWR.n1546 VGND 0.021519f
C6141 VDPWR.n1547 VGND 0.030925f
C6142 VDPWR.n1548 VGND 0.021519f
C6143 VDPWR.n1549 VGND 0.014025f
C6144 VDPWR.n1550 VGND 0.051783f
C6145 VDPWR.n1551 VGND 0.093119f
C6146 VDPWR.n1552 VGND 0.014025f
C6147 VDPWR.n1553 VGND 0.021519f
C6148 VDPWR.n1554 VGND 0.030925f
C6149 VDPWR.n1555 VGND 0.021519f
C6150 VDPWR.n1556 VGND 0.014025f
C6151 VDPWR.n1557 VGND 0.051783f
C6152 VDPWR.n1558 VGND 0.093119f
C6153 VDPWR.n1559 VGND 0.014025f
C6154 VDPWR.n1560 VGND 0.021519f
C6155 VDPWR.n1561 VGND 0.030925f
C6156 VDPWR.n1562 VGND 0.041191f
C6157 VDPWR.n1563 VGND 0.014025f
C6158 VDPWR.n1564 VGND 0.048444f
C6159 VDPWR.n1565 VGND 0.958126f
C6160 VDPWR.n1566 VGND 21.3883f
C6161 VDPWR.n1567 VGND 5.62448f
C6162 VDPWR.n1568 VGND 5.97167f
C6163 VDPWR.n1569 VGND 0.196532f
C6164 VDPWR.n1570 VGND 0.062518f
C6165 VDPWR.n1571 VGND 0.019706f
C6166 VDPWR.n1572 VGND 0.161177f
C6167 VDPWR.n1573 VGND 0.032123f
C6168 VDPWR.n1574 VGND 0.0501f
C6169 VDPWR.n1575 VGND 0.081439f
C6170 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 VGND 0.060722f
C6171 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 VGND 0.060722f
C6172 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 VGND 0.070899f
C6173 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 VGND 0.060722f
C6174 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 VGND 0.060722f
C6175 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 VGND 0.070523f
C6176 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 VGND 0.632153f
C6177 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 VGND 0.059856f
C6178 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 VGND 0.019094f
C6179 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 VGND 0.041709f
C6180 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 VGND 0.059856f
C6181 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 VGND 0.019094f
C6182 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 VGND 0.04198f
C6183 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 VGND 0.013454f
C6184 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 VGND 0.059856f
C6185 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 VGND 0.019094f
C6186 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 VGND 0.04198f
C6187 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 VGND 0.059856f
C6188 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 VGND 0.019094f
C6189 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 VGND 0.041709f
C6190 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 VGND 0.013307f
C6191 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 VGND 0.351257f
C6192 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 VGND 0.047903f
C6193 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 VGND 0.144997f
C6194 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 VGND 0.368007f
C6195 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 VGND 0.013091f
C6196 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 VGND 0.013091f
C6197 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 VGND 0.030662f
C6198 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 VGND 0.039272f
C6199 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 VGND 0.039272f
C6200 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 VGND 0.080004f
C6201 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 VGND 0.332866f
C6202 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 VGND 0.180864f
C6203 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 VGND 0.144997f
C6204 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 VGND 0.240639f
C6205 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 VGND 0.045973f
C6206 tdc_0.vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 VGND 0.156775f
.ends

